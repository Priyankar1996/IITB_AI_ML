-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_Block0_start_973_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1050_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1217_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_ack_0 : boolean;
  signal type_cast_733_inst_req_1 : boolean;
  signal type_cast_733_inst_ack_1 : boolean;
  signal type_cast_715_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1050_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_req_1 : boolean;
  signal type_cast_1035_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1214_inst_req_0 : boolean;
  signal type_cast_472_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1021_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_711_inst_req_0 : boolean;
  signal type_cast_526_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1015_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1277_inst_ack_1 : boolean;
  signal type_cast_733_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_747_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_540_inst_ack_1 : boolean;
  signal type_cast_526_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_540_inst_req_1 : boolean;
  signal type_cast_490_inst_ack_0 : boolean;
  signal type_cast_490_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_540_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_540_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_961_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal WPIPE_Block0_start_961_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal type_cast_715_inst_req_1 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_967_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_522_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_639_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_639_inst_req_1 : boolean;
  signal type_cast_51_inst_req_0 : boolean;
  signal type_cast_51_inst_ack_0 : boolean;
  signal type_cast_51_inst_req_1 : boolean;
  signal type_cast_51_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_988_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1003_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 : boolean;
  signal type_cast_526_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 : boolean;
  signal type_cast_1035_inst_req_1 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal type_cast_643_inst_ack_1 : boolean;
  signal type_cast_526_inst_req_0 : boolean;
  signal type_cast_593_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1003_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1027_inst_req_1 : boolean;
  signal type_cast_593_inst_req_1 : boolean;
  signal WPIPE_Block0_start_949_inst_req_0 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1027_inst_ack_1 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal array_obj_ref_622_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_967_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_639_inst_ack_0 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal type_cast_643_inst_req_1 : boolean;
  signal array_obj_ref_622_index_offset_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 : boolean;
  signal type_cast_715_inst_ack_0 : boolean;
  signal type_cast_679_inst_ack_1 : boolean;
  signal type_cast_679_inst_req_1 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_639_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_626_inst_ack_1 : boolean;
  signal type_cast_101_inst_req_0 : boolean;
  signal WPIPE_Block0_start_970_inst_req_0 : boolean;
  signal type_cast_101_inst_ack_0 : boolean;
  signal type_cast_101_inst_req_1 : boolean;
  signal type_cast_101_inst_ack_1 : boolean;
  signal array_obj_ref_622_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_657_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_522_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 : boolean;
  signal type_cast_679_inst_ack_0 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_626_inst_req_1 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_973_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_1 : boolean;
  signal WPIPE_Block1_start_988_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_522_inst_req_1 : boolean;
  signal array_obj_ref_622_index_offset_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_657_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 : boolean;
  signal type_cast_679_inst_req_0 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_0 : boolean;
  signal type_cast_643_inst_ack_0 : boolean;
  signal addr_of_623_final_reg_ack_0 : boolean;
  signal WPIPE_Block0_start_949_inst_req_1 : boolean;
  signal if_stmt_350_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1003_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_486_inst_req_0 : boolean;
  signal if_stmt_350_branch_ack_1 : boolean;
  signal if_stmt_350_branch_ack_0 : boolean;
  signal type_cast_138_inst_req_0 : boolean;
  signal type_cast_138_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_626_inst_ack_0 : boolean;
  signal type_cast_138_inst_req_1 : boolean;
  signal type_cast_138_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_522_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_1 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_991_inst_req_0 : boolean;
  signal type_cast_151_inst_req_0 : boolean;
  signal type_cast_151_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_626_inst_req_0 : boolean;
  signal type_cast_151_inst_req_1 : boolean;
  signal type_cast_151_inst_ack_1 : boolean;
  signal type_cast_697_inst_ack_1 : boolean;
  signal type_cast_643_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_729_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_949_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_657_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_657_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 : boolean;
  signal type_cast_163_inst_req_0 : boolean;
  signal type_cast_163_inst_ack_0 : boolean;
  signal type_cast_163_inst_req_1 : boolean;
  signal type_cast_163_inst_ack_1 : boolean;
  signal type_cast_697_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_729_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 : boolean;
  signal type_cast_715_inst_req_0 : boolean;
  signal type_cast_176_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1243_inst_req_0 : boolean;
  signal type_cast_176_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1015_inst_req_0 : boolean;
  signal type_cast_176_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 : boolean;
  signal type_cast_508_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1024_inst_req_1 : boolean;
  signal WPIPE_Block1_start_991_inst_ack_1 : boolean;
  signal type_cast_188_inst_req_0 : boolean;
  signal type_cast_188_inst_ack_0 : boolean;
  signal type_cast_188_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1015_inst_ack_0 : boolean;
  signal type_cast_188_inst_ack_1 : boolean;
  signal type_cast_508_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1217_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1024_inst_ack_1 : boolean;
  signal type_cast_201_inst_req_0 : boolean;
  signal type_cast_201_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_961_inst_ack_1 : boolean;
  signal type_cast_201_inst_req_1 : boolean;
  signal ptr_deref_552_store_0_ack_1 : boolean;
  signal type_cast_201_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_967_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_729_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1243_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_257_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_257_inst_ack_0 : boolean;
  signal type_cast_508_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_257_inst_req_1 : boolean;
  signal ptr_deref_552_store_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_257_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_675_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_675_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_260_inst_req_0 : boolean;
  signal WPIPE_Block0_start_970_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_260_inst_ack_0 : boolean;
  signal type_cast_508_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_260_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_260_inst_ack_1 : boolean;
  signal type_cast_1035_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_263_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1003_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_675_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_675_inst_req_0 : boolean;
  signal type_cast_630_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_266_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_266_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_266_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_266_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_711_inst_ack_1 : boolean;
  signal type_cast_630_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_269_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_269_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_269_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_269_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_711_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_994_inst_req_0 : boolean;
  signal WPIPE_Block1_start_994_inst_ack_0 : boolean;
  signal type_cast_273_inst_req_0 : boolean;
  signal type_cast_273_inst_ack_0 : boolean;
  signal type_cast_273_inst_req_1 : boolean;
  signal type_cast_273_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_729_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_req_1 : boolean;
  signal ptr_deref_552_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_ack_1 : boolean;
  signal type_cast_630_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_req_1 : boolean;
  signal if_stmt_566_branch_ack_0 : boolean;
  signal type_cast_286_inst_req_0 : boolean;
  signal type_cast_286_inst_ack_0 : boolean;
  signal type_cast_286_inst_req_1 : boolean;
  signal ptr_deref_552_store_0_req_0 : boolean;
  signal type_cast_286_inst_ack_1 : boolean;
  signal type_cast_697_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_967_inst_req_0 : boolean;
  signal WPIPE_Block0_start_949_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_504_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_957_inst_req_1 : boolean;
  signal type_cast_630_inst_req_0 : boolean;
  signal type_cast_298_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_504_inst_req_1 : boolean;
  signal type_cast_298_inst_ack_0 : boolean;
  signal type_cast_298_inst_req_1 : boolean;
  signal type_cast_298_inst_ack_1 : boolean;
  signal type_cast_697_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_req_0 : boolean;
  signal WPIPE_Block0_start_970_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_957_inst_ack_1 : boolean;
  signal if_stmt_566_branch_ack_1 : boolean;
  signal type_cast_544_inst_ack_1 : boolean;
  signal type_cast_311_inst_req_0 : boolean;
  signal type_cast_311_inst_ack_0 : boolean;
  signal type_cast_311_inst_req_1 : boolean;
  signal type_cast_311_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_504_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_319_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_319_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_504_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_319_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_319_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_711_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1053_inst_req_0 : boolean;
  signal type_cast_661_inst_ack_1 : boolean;
  signal type_cast_661_inst_req_1 : boolean;
  signal type_cast_544_inst_req_1 : boolean;
  signal type_cast_323_inst_req_0 : boolean;
  signal type_cast_323_inst_ack_0 : boolean;
  signal type_cast_323_inst_req_1 : boolean;
  signal type_cast_323_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1187_inst_req_1 : boolean;
  signal WPIPE_Block1_start_991_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_332_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_332_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_332_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_332_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_991_inst_ack_0 : boolean;
  signal type_cast_336_inst_req_0 : boolean;
  signal type_cast_336_inst_ack_0 : boolean;
  signal type_cast_336_inst_req_1 : boolean;
  signal type_cast_336_inst_ack_1 : boolean;
  signal type_cast_661_inst_ack_0 : boolean;
  signal type_cast_661_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1255_inst_ack_0 : boolean;
  signal addr_of_623_final_reg_ack_1 : boolean;
  signal if_stmt_365_branch_req_0 : boolean;
  signal if_stmt_365_branch_ack_1 : boolean;
  signal if_stmt_365_branch_ack_0 : boolean;
  signal addr_of_623_final_reg_req_1 : boolean;
  signal type_cast_386_inst_req_0 : boolean;
  signal type_cast_386_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1214_inst_ack_1 : boolean;
  signal type_cast_386_inst_req_1 : boolean;
  signal type_cast_386_inst_ack_1 : boolean;
  signal type_cast_733_inst_req_0 : boolean;
  signal type_cast_544_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_994_inst_req_1 : boolean;
  signal addr_of_623_final_reg_req_0 : boolean;
  signal type_cast_544_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_994_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_693_inst_req_0 : boolean;
  signal array_obj_ref_415_index_offset_req_0 : boolean;
  signal array_obj_ref_415_index_offset_ack_0 : boolean;
  signal array_obj_ref_415_index_offset_req_1 : boolean;
  signal array_obj_ref_415_index_offset_ack_1 : boolean;
  signal WPIPE_Block3_start_1264_inst_ack_1 : boolean;
  signal addr_of_416_final_reg_req_0 : boolean;
  signal addr_of_416_final_reg_ack_0 : boolean;
  signal addr_of_416_final_reg_req_1 : boolean;
  signal addr_of_416_final_reg_ack_1 : boolean;
  signal if_stmt_566_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_419_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_419_inst_ack_0 : boolean;
  signal type_cast_490_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_419_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_419_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1053_inst_ack_0 : boolean;
  signal type_cast_423_inst_req_0 : boolean;
  signal type_cast_423_inst_ack_0 : boolean;
  signal type_cast_423_inst_req_1 : boolean;
  signal type_cast_490_inst_req_1 : boolean;
  signal type_cast_423_inst_ack_1 : boolean;
  signal type_cast_472_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_976_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_432_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_432_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_970_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_432_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_432_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_961_inst_req_1 : boolean;
  signal type_cast_436_inst_req_0 : boolean;
  signal type_cast_436_inst_ack_0 : boolean;
  signal type_cast_436_inst_req_1 : boolean;
  signal type_cast_436_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_450_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_450_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_450_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_450_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_997_inst_req_0 : boolean;
  signal type_cast_454_inst_req_0 : boolean;
  signal type_cast_454_inst_ack_0 : boolean;
  signal type_cast_454_inst_req_1 : boolean;
  signal type_cast_454_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_468_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_468_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_468_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_468_inst_ack_1 : boolean;
  signal type_cast_472_inst_req_0 : boolean;
  signal type_cast_472_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_957_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_988_inst_ack_0 : boolean;
  signal type_cast_751_inst_req_0 : boolean;
  signal type_cast_751_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1217_inst_ack_1 : boolean;
  signal type_cast_751_inst_req_1 : boolean;
  signal type_cast_751_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1059_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1018_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1018_inst_req_1 : boolean;
  signal WPIPE_Block1_start_988_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1021_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1027_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1243_inst_req_1 : boolean;
  signal WPIPE_Block0_start_973_inst_ack_0 : boolean;
  signal ptr_deref_759_store_0_req_0 : boolean;
  signal ptr_deref_759_store_0_ack_0 : boolean;
  signal ptr_deref_759_store_0_req_1 : boolean;
  signal ptr_deref_759_store_0_ack_1 : boolean;
  signal WPIPE_Block1_start_1059_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1268_inst_req_0 : boolean;
  signal WPIPE_Block0_start_957_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1027_inst_req_0 : boolean;
  signal if_stmt_773_branch_req_0 : boolean;
  signal type_cast_1035_inst_req_0 : boolean;
  signal if_stmt_773_branch_ack_1 : boolean;
  signal if_stmt_773_branch_ack_0 : boolean;
  signal WPIPE_Block0_start_973_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1000_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1000_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_ack_1 : boolean;
  signal if_stmt_798_branch_req_0 : boolean;
  signal WPIPE_Block1_start_985_inst_ack_1 : boolean;
  signal if_stmt_798_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1000_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_1 : boolean;
  signal if_stmt_798_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1056_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1000_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1018_inst_ack_0 : boolean;
  signal type_cast_825_inst_req_0 : boolean;
  signal type_cast_825_inst_ack_0 : boolean;
  signal type_cast_825_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1199_inst_req_0 : boolean;
  signal type_cast_825_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1021_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1024_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_985_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1018_inst_req_0 : boolean;
  signal WPIPE_Block0_start_953_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1053_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1053_inst_req_1 : boolean;
  signal WPIPE_Block1_start_985_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1021_inst_req_0 : boolean;
  signal array_obj_ref_854_index_offset_req_0 : boolean;
  signal WPIPE_Block1_start_1012_inst_ack_1 : boolean;
  signal array_obj_ref_854_index_offset_ack_0 : boolean;
  signal array_obj_ref_854_index_offset_req_1 : boolean;
  signal array_obj_ref_854_index_offset_ack_1 : boolean;
  signal WPIPE_Block1_start_1024_inst_req_0 : boolean;
  signal WPIPE_Block1_start_985_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1012_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1243_inst_ack_1 : boolean;
  signal addr_of_855_final_reg_req_0 : boolean;
  signal addr_of_855_final_reg_ack_0 : boolean;
  signal addr_of_855_final_reg_req_1 : boolean;
  signal addr_of_855_final_reg_ack_1 : boolean;
  signal WPIPE_Block3_start_1252_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1255_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1255_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1012_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1196_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1012_inst_req_0 : boolean;
  signal ptr_deref_858_store_0_req_0 : boolean;
  signal ptr_deref_858_store_0_ack_0 : boolean;
  signal ptr_deref_858_store_0_req_1 : boolean;
  signal ptr_deref_858_store_0_ack_1 : boolean;
  signal WPIPE_Block3_start_1261_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_982_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_997_inst_ack_1 : boolean;
  signal if_stmt_873_branch_req_0 : boolean;
  signal WPIPE_Block3_start_1214_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_982_inst_req_1 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_997_inst_req_1 : boolean;
  signal WPIPE_Block0_start_953_inst_req_0 : boolean;
  signal if_stmt_873_branch_ack_1 : boolean;
  signal if_stmt_873_branch_ack_0 : boolean;
  signal call_stmt_884_call_req_0 : boolean;
  signal call_stmt_884_call_ack_0 : boolean;
  signal call_stmt_884_call_req_1 : boolean;
  signal call_stmt_884_call_ack_1 : boolean;
  signal type_cast_889_inst_req_0 : boolean;
  signal type_cast_889_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_997_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1255_inst_req_0 : boolean;
  signal type_cast_889_inst_req_1 : boolean;
  signal type_cast_889_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_891_inst_req_0 : boolean;
  signal WPIPE_Block0_start_891_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_891_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1009_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_891_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_894_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1009_inst_req_1 : boolean;
  signal WPIPE_Block0_start_894_inst_ack_0 : boolean;
  signal type_cast_1048_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_894_inst_req_1 : boolean;
  signal WPIPE_Block0_start_894_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1264_inst_req_1 : boolean;
  signal WPIPE_Block1_start_982_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_897_inst_req_0 : boolean;
  signal WPIPE_Block0_start_897_inst_ack_0 : boolean;
  signal type_cast_1048_inst_req_1 : boolean;
  signal WPIPE_Block0_start_897_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1009_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_897_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1214_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_982_inst_req_0 : boolean;
  signal WPIPE_Block0_start_900_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1009_inst_req_0 : boolean;
  signal WPIPE_Block0_start_900_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_900_inst_req_1 : boolean;
  signal WPIPE_Block0_start_900_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1050_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_req_0 : boolean;
  signal WPIPE_Block0_start_903_inst_req_0 : boolean;
  signal WPIPE_Block0_start_903_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_964_inst_ack_1 : boolean;
  signal type_cast_1048_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_903_inst_req_1 : boolean;
  signal WPIPE_Block0_start_903_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1050_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1187_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1217_inst_req_0 : boolean;
  signal WPIPE_Block0_start_906_inst_req_0 : boolean;
  signal WPIPE_Block0_start_906_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_964_inst_req_1 : boolean;
  signal type_cast_1048_inst_req_0 : boolean;
  signal WPIPE_Block0_start_906_inst_req_1 : boolean;
  signal WPIPE_Block0_start_906_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1015_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_909_inst_req_0 : boolean;
  signal WPIPE_Block0_start_909_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_909_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1006_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_909_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1030_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_912_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1006_inst_req_1 : boolean;
  signal WPIPE_Block0_start_912_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_912_inst_req_1 : boolean;
  signal WPIPE_Block0_start_912_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1264_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1030_inst_req_1 : boolean;
  signal WPIPE_Block1_start_979_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_979_inst_req_1 : boolean;
  signal WPIPE_Block0_start_915_inst_req_0 : boolean;
  signal WPIPE_Block0_start_915_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_915_inst_req_1 : boolean;
  signal WPIPE_Block0_start_915_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_964_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1030_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_979_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_979_inst_req_0 : boolean;
  signal WPIPE_Block0_start_918_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1006_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_918_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_964_inst_req_0 : boolean;
  signal WPIPE_Block0_start_918_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1006_inst_req_0 : boolean;
  signal WPIPE_Block0_start_918_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1030_inst_req_0 : boolean;
  signal WPIPE_Block0_start_921_inst_req_0 : boolean;
  signal WPIPE_Block0_start_921_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_921_inst_req_1 : boolean;
  signal WPIPE_Block0_start_921_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1277_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1268_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_924_inst_req_0 : boolean;
  signal WPIPE_Block0_start_924_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_924_inst_req_1 : boolean;
  signal WPIPE_Block0_start_924_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1196_inst_req_1 : boolean;
  signal WPIPE_Block0_start_976_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_976_inst_req_1 : boolean;
  signal WPIPE_Block0_start_927_inst_req_0 : boolean;
  signal WPIPE_Block0_start_927_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_927_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1199_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_927_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1187_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_930_inst_req_0 : boolean;
  signal WPIPE_Block0_start_930_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1277_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_930_inst_req_1 : boolean;
  signal WPIPE_Block0_start_930_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1268_inst_req_1 : boolean;
  signal WPIPE_Block0_start_933_inst_req_0 : boolean;
  signal WPIPE_Block0_start_933_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_933_inst_req_1 : boolean;
  signal WPIPE_Block0_start_933_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1199_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1199_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_936_inst_req_0 : boolean;
  signal WPIPE_Block0_start_936_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_936_inst_req_1 : boolean;
  signal WPIPE_Block0_start_936_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1277_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1246_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1246_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_939_inst_req_0 : boolean;
  signal WPIPE_Block0_start_939_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_939_inst_req_1 : boolean;
  signal WPIPE_Block0_start_939_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_942_inst_req_0 : boolean;
  signal WPIPE_Block0_start_942_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_942_inst_req_1 : boolean;
  signal WPIPE_Block0_start_942_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_945_inst_req_0 : boolean;
  signal WPIPE_Block0_start_945_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_945_inst_req_1 : boolean;
  signal WPIPE_Block0_start_945_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1059_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1059_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1160_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1252_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1062_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1240_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1062_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1062_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1240_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1062_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1065_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1065_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1065_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1065_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1211_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1211_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1068_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1240_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1068_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1196_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1068_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1240_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1068_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1274_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1252_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1261_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1071_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1071_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1196_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1071_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1071_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1274_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1252_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1074_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1074_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1074_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1074_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1211_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1077_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1077_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1077_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1077_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1211_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1261_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1080_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1080_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1080_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1080_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1274_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1261_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1083_inst_req_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1083_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1083_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1083_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1274_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1086_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1086_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1086_inst_req_1 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1086_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1089_inst_req_0 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1089_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1089_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1089_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1092_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1092_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1193_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1092_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1092_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1249_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1095_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1095_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1193_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1095_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1095_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1249_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1098_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1098_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1098_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1226_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1098_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1208_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1101_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1101_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1101_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1226_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1101_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1208_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1258_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1104_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1104_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1104_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1104_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1249_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1258_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1107_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1226_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1107_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1193_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1107_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1226_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1107_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1249_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1110_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1110_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1193_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1110_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1110_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1208_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1113_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1113_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1271_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1208_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1258_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1116_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1116_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1271_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1258_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1223_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1223_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1271_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1223_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1223_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1271_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1128_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1205_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1131_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1131_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1190_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1131_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1131_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1205_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1246_inst_ack_1 : boolean;
  signal type_cast_1143_inst_req_0 : boolean;
  signal type_cast_1143_inst_ack_0 : boolean;
  signal type_cast_1143_inst_req_1 : boolean;
  signal type_cast_1143_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1190_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1246_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1205_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1145_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1220_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1145_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1145_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1220_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1145_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1190_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1205_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1148_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1148_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1190_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1148_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1148_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1151_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1220_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1151_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1151_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1220_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1151_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1202_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1264_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1202_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1154_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1154_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1154_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1154_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1202_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1202_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1157_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1157_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1157_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1157_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1187_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1268_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1160_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1160_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1160_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1163_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1163_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1163_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1163_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1166_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1166_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1166_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1166_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1169_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1169_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1169_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1169_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1172_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1172_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1172_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1172_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_1 : boolean;
  signal call_stmt_1281_call_req_0 : boolean;
  signal call_stmt_1281_call_ack_0 : boolean;
  signal call_stmt_1281_call_req_1 : boolean;
  signal call_stmt_1281_call_ack_1 : boolean;
  signal type_cast_1285_inst_req_0 : boolean;
  signal type_cast_1285_inst_ack_0 : boolean;
  signal type_cast_1285_inst_req_1 : boolean;
  signal type_cast_1285_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1292_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1292_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1292_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1292_inst_ack_1 : boolean;
  signal phi_stmt_1340_req_0 : boolean;
  signal if_stmt_1296_branch_req_0 : boolean;
  signal if_stmt_1296_branch_ack_1 : boolean;
  signal if_stmt_1296_branch_ack_0 : boolean;
  signal type_cast_1323_inst_req_0 : boolean;
  signal type_cast_1323_inst_ack_0 : boolean;
  signal type_cast_1323_inst_req_1 : boolean;
  signal type_cast_1323_inst_ack_1 : boolean;
  signal array_obj_ref_1352_index_offset_req_0 : boolean;
  signal array_obj_ref_1352_index_offset_ack_0 : boolean;
  signal array_obj_ref_1352_index_offset_req_1 : boolean;
  signal array_obj_ref_1352_index_offset_ack_1 : boolean;
  signal addr_of_1353_final_reg_req_0 : boolean;
  signal addr_of_1353_final_reg_ack_0 : boolean;
  signal addr_of_1353_final_reg_req_1 : boolean;
  signal addr_of_1353_final_reg_ack_1 : boolean;
  signal ptr_deref_1357_load_0_req_0 : boolean;
  signal ptr_deref_1357_load_0_ack_0 : boolean;
  signal ptr_deref_1357_load_0_req_1 : boolean;
  signal ptr_deref_1357_load_0_ack_1 : boolean;
  signal phi_stmt_1340_ack_0 : boolean;
  signal type_cast_1361_inst_req_0 : boolean;
  signal type_cast_1361_inst_ack_0 : boolean;
  signal type_cast_1361_inst_req_1 : boolean;
  signal type_cast_1361_inst_ack_1 : boolean;
  signal type_cast_1371_inst_req_0 : boolean;
  signal type_cast_1371_inst_ack_0 : boolean;
  signal type_cast_1371_inst_req_1 : boolean;
  signal type_cast_1371_inst_ack_1 : boolean;
  signal phi_stmt_1340_req_1 : boolean;
  signal type_cast_1346_inst_ack_1 : boolean;
  signal type_cast_1381_inst_req_0 : boolean;
  signal type_cast_1381_inst_ack_0 : boolean;
  signal type_cast_1381_inst_req_1 : boolean;
  signal type_cast_1381_inst_ack_1 : boolean;
  signal type_cast_1346_inst_req_1 : boolean;
  signal type_cast_1391_inst_req_0 : boolean;
  signal type_cast_1391_inst_ack_0 : boolean;
  signal type_cast_1391_inst_req_1 : boolean;
  signal type_cast_1391_inst_ack_1 : boolean;
  signal type_cast_1346_inst_ack_0 : boolean;
  signal type_cast_1401_inst_req_0 : boolean;
  signal type_cast_1401_inst_ack_0 : boolean;
  signal type_cast_1346_inst_req_0 : boolean;
  signal type_cast_1401_inst_req_1 : boolean;
  signal type_cast_1401_inst_ack_1 : boolean;
  signal type_cast_1411_inst_req_0 : boolean;
  signal type_cast_1411_inst_ack_0 : boolean;
  signal type_cast_1411_inst_req_1 : boolean;
  signal type_cast_1411_inst_ack_1 : boolean;
  signal type_cast_1421_inst_req_0 : boolean;
  signal type_cast_1421_inst_ack_0 : boolean;
  signal type_cast_1421_inst_req_1 : boolean;
  signal type_cast_1421_inst_ack_1 : boolean;
  signal type_cast_1431_inst_req_0 : boolean;
  signal type_cast_1431_inst_ack_0 : boolean;
  signal type_cast_1431_inst_req_1 : boolean;
  signal type_cast_1431_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1433_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1433_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1433_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1433_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1436_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1436_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1436_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1436_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1439_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1439_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1439_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1439_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1 : boolean;
  signal if_stmt_1468_branch_req_0 : boolean;
  signal if_stmt_1468_branch_ack_1 : boolean;
  signal if_stmt_1468_branch_ack_0 : boolean;
  signal phi_stmt_403_req_0 : boolean;
  signal type_cast_409_inst_req_0 : boolean;
  signal type_cast_409_inst_ack_0 : boolean;
  signal type_cast_409_inst_req_1 : boolean;
  signal type_cast_409_inst_ack_1 : boolean;
  signal phi_stmt_403_req_1 : boolean;
  signal phi_stmt_403_ack_0 : boolean;
  signal phi_stmt_610_req_0 : boolean;
  signal type_cast_616_inst_req_0 : boolean;
  signal type_cast_616_inst_ack_0 : boolean;
  signal type_cast_616_inst_req_1 : boolean;
  signal type_cast_616_inst_ack_1 : boolean;
  signal phi_stmt_610_req_1 : boolean;
  signal phi_stmt_610_ack_0 : boolean;
  signal phi_stmt_842_req_0 : boolean;
  signal type_cast_848_inst_req_0 : boolean;
  signal type_cast_848_inst_ack_0 : boolean;
  signal type_cast_848_inst_req_1 : boolean;
  signal type_cast_848_inst_ack_1 : boolean;
  signal phi_stmt_842_req_1 : boolean;
  signal phi_stmt_842_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(535 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(535);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	80 
    -- CP-element group 0: 	72 
    -- CP-element group 0: 	84 
    -- CP-element group 0: 	88 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (68) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_Update/cr
      -- 
    rr_133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_51_inst_req_1); -- 
    cr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_63_inst_req_1); -- 
    cr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_76_inst_req_1); -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_88_inst_req_1); -- 
    cr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_101_inst_req_1); -- 
    cr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_113_inst_req_1); -- 
    cr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_126_inst_req_1); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_138_inst_req_1); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_151_inst_req_1); -- 
    cr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_163_inst_req_1); -- 
    cr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_176_inst_req_1); -- 
    cr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_188_inst_req_1); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_201_inst_req_1); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_273_inst_req_1); -- 
    cr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_286_inst_req_1); -- 
    cr_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_298_inst_req_1); -- 
    cr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_311_inst_req_1); -- 
    cr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_323_inst_req_1); -- 
    cr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_336_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_Sample/rr
      -- 
    ca_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_Sample/ra
      -- 
    ra_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	89 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_38_Update/ca
      -- 
    ca_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_update_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_Update/cr
      -- 
    ra_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_47_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_Sample/rr
      -- 
    ca_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_51_inst_req_0); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_Sample/ra
      -- 
    ra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	89 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_51_Update/ca
      -- 
    ca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_update_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_Update/cr
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_59_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_Sample/rr
      -- 
    ca_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_63_inst_req_0); -- 
    rr_217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_Sample/ra
      -- 
    ra_204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	89 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_63_Update/ca
      -- 
    ca_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_update_start_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_Update/cr
      -- 
    ra_218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_72_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_Sample/rr
      -- 
    ca_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_76_inst_req_0); -- 
    rr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_Sample/ra
      -- 
    ra_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	89 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_76_Update/ca
      -- 
    ca_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_update_start_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_Update/cr
      -- 
    ra_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_84_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_Sample/rr
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_88_inst_req_0); -- 
    rr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_Sample/ra
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	89 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_88_Update/ca
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_update_start_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_Update/cr
      -- 
    ra_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_97_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_Sample/rr
      -- 
    ca_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_101_inst_req_0); -- 
    rr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_Sample/ra
      -- 
    ra_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	89 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_101_Update/ca
      -- 
    ca_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_update_start_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_Update/cr
      -- 
    ra_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_109_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_Sample/rr
      -- 
    ca_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_113_inst_req_0); -- 
    rr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_Sample/ra
      -- 
    ra_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	89 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_113_Update/ca
      -- 
    ca_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_update_start_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_Update/cr
      -- 
    ra_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_122_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_Sample/$entry
      -- 
    ca_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_126_inst_req_0); -- 
    rr_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_Sample/ra
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	89 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_126_Update/ca
      -- 
    ca_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_update_start_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_Sample/$exit
      -- 
    ra_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_134_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_Sample/rr
      -- 
    ca_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_138_inst_req_0); -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_Sample/ra
      -- 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	89 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_138_Update/ca
      -- 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_update_start_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_Update/cr
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_147_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_Sample/rr
      -- 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_0); -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_151_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	89 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_151_Update/ca
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_update_start_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_Update/cr
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_159_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_Sample/rr
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_0); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_163_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_Sample/ra
      -- 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	89 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_163_Update/ca
      -- 
    ca_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_update_start_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_Update/cr
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_172_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_Sample/rr
      -- 
    ca_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_176_inst_req_0); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_Sample/ra
      -- 
    ra_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	89 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_176_Update/ca
      -- 
    ca_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_update_start_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_Update/cr
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_184_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_Sample/rr
      -- 
    ca_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_0); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_188_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_Sample/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	89 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_188_Update/ca
      -- 
    ca_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_update_start_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_Update/cr
      -- 
    ra_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_197_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_Sample/rr
      -- 
    ca_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_201_inst_req_0); -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_257_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_Sample/ra
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	89 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_201_Update/ca
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_update_start_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_Update/cr
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_257_inst_ack_0, ack => convTranspose_CP_39_elements(57)); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => RPIPE_ConvTranspose_input_pipe_257_inst_req_1); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_257_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_Sample/rr
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_257_inst_ack_1, ack => convTranspose_CP_39_elements(58)); -- 
    rr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(58), ack => RPIPE_ConvTranspose_input_pipe_260_inst_req_0); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_update_start_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_Sample/ra
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_Update/cr
      -- 
    ra_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_260_inst_ack_0, ack => convTranspose_CP_39_elements(59)); -- 
    cr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(59), ack => RPIPE_ConvTranspose_input_pipe_260_inst_req_1); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_260_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_Sample/rr
      -- 
    ca_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_260_inst_ack_1, ack => convTranspose_CP_39_elements(60)); -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(60), ack => RPIPE_ConvTranspose_input_pipe_263_inst_req_0); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_update_start_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_Update/cr
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_263_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(61), ack => RPIPE_ConvTranspose_input_pipe_263_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_263_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_Sample/rr
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_263_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    rr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(62), ack => RPIPE_ConvTranspose_input_pipe_266_inst_req_0); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_update_start_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_Update/cr
      -- 
    ra_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_266_inst_ack_0, ack => convTranspose_CP_39_elements(63)); -- 
    cr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(63), ack => RPIPE_ConvTranspose_input_pipe_266_inst_req_1); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_266_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_Sample/rr
      -- 
    ca_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_266_inst_ack_1, ack => convTranspose_CP_39_elements(64)); -- 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(64), ack => RPIPE_ConvTranspose_input_pipe_269_inst_req_0); -- 
    -- CP-element group 65:  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_update_start_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_Update/cr
      -- 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_269_inst_ack_0, ack => convTranspose_CP_39_elements(65)); -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(65), ack => RPIPE_ConvTranspose_input_pipe_269_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	69 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_269_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_Sample/rr
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_269_inst_ack_1, ack => convTranspose_CP_39_elements(66)); -- 
    rr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => RPIPE_ConvTranspose_input_pipe_282_inst_req_0); -- 
    rr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_273_inst_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_Sample/ra
      -- 
    ra_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	89 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_273_Update/ca
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	66 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_update_start_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_Update/cr
      -- 
    ra_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_282_inst_ack_0, ack => convTranspose_CP_39_elements(69)); -- 
    cr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => RPIPE_ConvTranspose_input_pipe_282_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	73 
    -- CP-element group 70:  members (9) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_282_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_Sample/rr
      -- 
    ca_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_282_inst_ack_1, ack => convTranspose_CP_39_elements(70)); -- 
    rr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(70), ack => type_cast_286_inst_req_0); -- 
    rr_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(70), ack => RPIPE_ConvTranspose_input_pipe_294_inst_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_Sample/ra
      -- 
    ra_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_286_inst_ack_0, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	0 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	89 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_286_Update/ca
      -- 
    ca_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_286_inst_ack_1, ack => convTranspose_CP_39_elements(72)); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	70 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_Update/cr
      -- 
    ra_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_294_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    cr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(73), ack => RPIPE_ConvTranspose_input_pipe_294_inst_req_1); -- 
    -- CP-element group 74:  fork  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	77 
    -- CP-element group 74:  members (9) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_294_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_Sample/rr
      -- 
    ca_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_294_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    rr_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(74), ack => RPIPE_ConvTranspose_input_pipe_307_inst_req_0); -- 
    rr_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(74), ack => type_cast_298_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_Sample/ra
      -- 
    ra_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_298_inst_ack_0, ack => convTranspose_CP_39_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	89 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_298_Update/ca
      -- 
    ca_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_298_inst_ack_1, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	74 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_Update/cr
      -- 
    ra_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_307_inst_ack_0, ack => convTranspose_CP_39_elements(77)); -- 
    cr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(77), ack => RPIPE_ConvTranspose_input_pipe_307_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	81 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_307_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_Sample/rr
      -- 
    ca_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_307_inst_ack_1, ack => convTranspose_CP_39_elements(78)); -- 
    rr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => type_cast_311_inst_req_0); -- 
    rr_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_319_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_Sample/ra
      -- 
    ra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_0, ack => convTranspose_CP_39_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	0 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	89 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_311_Update/ca
      -- 
    ca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_1, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	78 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_update_start_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_Update/cr
      -- 
    ra_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_319_inst_ack_0, ack => convTranspose_CP_39_elements(81)); -- 
    cr_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(81), ack => RPIPE_ConvTranspose_input_pipe_319_inst_req_1); -- 
    -- CP-element group 82:  fork  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_319_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_Sample/rr
      -- 
    ca_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_319_inst_ack_1, ack => convTranspose_CP_39_elements(82)); -- 
    rr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => type_cast_323_inst_req_0); -- 
    rr_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_332_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_Sample/ra
      -- 
    ra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_323_inst_ack_0, ack => convTranspose_CP_39_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	0 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	89 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_323_Update/ca
      -- 
    ca_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_323_inst_ack_1, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	82 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_update_start_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_Sample/ra
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_Update/cr
      -- 
    ra_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_332_inst_ack_0, ack => convTranspose_CP_39_elements(85)); -- 
    cr_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(85), ack => RPIPE_ConvTranspose_input_pipe_332_inst_req_1); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/RPIPE_ConvTranspose_input_pipe_332_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_Sample/rr
      -- 
    ca_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_332_inst_ack_1, ack => convTranspose_CP_39_elements(86)); -- 
    rr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => type_cast_336_inst_req_0); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_Sample/ra
      -- 
    ra_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_336_inst_ack_0, ack => convTranspose_CP_39_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	0 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/type_cast_336_Update/ca
      -- 
    ca_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_336_inst_ack_1, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  branch  join  transition  place  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	44 
    -- CP-element group 89: 	68 
    -- CP-element group 89: 	40 
    -- CP-element group 89: 	52 
    -- CP-element group 89: 	48 
    -- CP-element group 89: 	56 
    -- CP-element group 89: 	76 
    -- CP-element group 89: 	80 
    -- CP-element group 89: 	72 
    -- CP-element group 89: 	84 
    -- CP-element group 89: 	88 
    -- CP-element group 89: 	4 
    -- CP-element group 89: 	8 
    -- CP-element group 89: 	12 
    -- CP-element group 89: 	16 
    -- CP-element group 89: 	20 
    -- CP-element group 89: 	24 
    -- CP-element group 89: 	28 
    -- CP-element group 89: 	32 
    -- CP-element group 89: 	36 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (10) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349__exit__
      -- CP-element group 89: 	 branch_block_stmt_32/if_stmt_350__entry__
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_349/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/if_stmt_350_dead_link/$entry
      -- CP-element group 89: 	 branch_block_stmt_32/if_stmt_350_eval_test/$entry
      -- CP-element group 89: 	 branch_block_stmt_32/if_stmt_350_eval_test/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/if_stmt_350_eval_test/branch_req
      -- CP-element group 89: 	 branch_block_stmt_32/R_cmp763_351_place
      -- CP-element group 89: 	 branch_block_stmt_32/if_stmt_350_if_link/$entry
      -- CP-element group 89: 	 branch_block_stmt_32/if_stmt_350_else_link/$entry
      -- 
    branch_req_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(89), ack => if_stmt_350_branch_req_0); -- 
    convTranspose_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 19) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1);
      constant place_markings: IntegerArray(0 to 19)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0);
      constant place_delays: IntegerArray(0 to 19) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 20); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(44) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(52) & convTranspose_CP_39_elements(48) & convTranspose_CP_39_elements(56) & convTranspose_CP_39_elements(76) & convTranspose_CP_39_elements(80) & convTranspose_CP_39_elements(72) & convTranspose_CP_39_elements(84) & convTranspose_CP_39_elements(88) & convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8) & convTranspose_CP_39_elements(12) & convTranspose_CP_39_elements(16) & convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(24) & convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(32) & convTranspose_CP_39_elements(36);
      gj_convTranspose_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 20, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90: 	95 
    -- CP-element group 90:  members (18) 
      -- CP-element group 90: 	 branch_block_stmt_32/merge_stmt_371__exit__
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400__entry__
      -- CP-element group 90: 	 branch_block_stmt_32/if_stmt_350_if_link/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/if_stmt_350_if_link/if_choice_transition
      -- CP-element group 90: 	 branch_block_stmt_32/entry_bbx_xnph765
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_update_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_Update/cr
      -- CP-element group 90: 	 branch_block_stmt_32/entry_bbx_xnph765_PhiReq/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/entry_bbx_xnph765_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/merge_stmt_371_PhiReqMerge
      -- CP-element group 90: 	 branch_block_stmt_32/merge_stmt_371_PhiAck/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/merge_stmt_371_PhiAck/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/merge_stmt_371_PhiAck/dummy
      -- 
    if_choice_transition_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_350_branch_ack_1, ack => convTranspose_CP_39_elements(90)); -- 
    rr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => type_cast_386_inst_req_0); -- 
    cr_798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => type_cast_386_inst_req_1); -- 
    -- CP-element group 91:  transition  place  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	508 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_32/if_stmt_350_else_link/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/if_stmt_350_else_link/else_choice_transition
      -- CP-element group 91: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader
      -- CP-element group 91: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_350_branch_ack_0, ack => convTranspose_CP_39_elements(91)); -- 
    -- CP-element group 92:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	508 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	138 
    -- CP-element group 92: 	139 
    -- CP-element group 92:  members (18) 
      -- CP-element group 92: 	 branch_block_stmt_32/merge_stmt_572__exit__
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607__entry__
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_update_start_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/$entry
      -- CP-element group 92: 	 branch_block_stmt_32/if_stmt_365_if_link/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/if_stmt_365_if_link/if_choice_transition
      -- CP-element group 92: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph761
      -- CP-element group 92: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph761_PhiReq/$entry
      -- CP-element group 92: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph761_PhiReq/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/merge_stmt_572_PhiReqMerge
      -- CP-element group 92: 	 branch_block_stmt_32/merge_stmt_572_PhiAck/$entry
      -- CP-element group 92: 	 branch_block_stmt_32/merge_stmt_572_PhiAck/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/merge_stmt_572_PhiAck/dummy
      -- 
    if_choice_transition_776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_365_branch_ack_1, ack => convTranspose_CP_39_elements(92)); -- 
    cr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(92), ack => type_cast_593_inst_req_1); -- 
    rr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(92), ack => type_cast_593_inst_req_0); -- 
    -- CP-element group 93:  transition  place  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	508 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	521 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_32/if_stmt_365_else_link/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/if_stmt_365_else_link/else_choice_transition
      -- CP-element group 93: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 93: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 93: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_365_branch_ack_0, ack => convTranspose_CP_39_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	90 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_Sample/ra
      -- 
    ra_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_386_inst_ack_0, ack => convTranspose_CP_39_elements(94)); -- 
    -- CP-element group 95:  transition  place  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	90 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	509 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400__exit__
      -- CP-element group 95: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_377_to_assign_stmt_400/type_cast_386_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody_PhiReq/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody_PhiReq/phi_stmt_403/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/$entry
      -- 
    ca_799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_386_inst_ack_1, ack => convTranspose_CP_39_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	514 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	135 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_sample_complete
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_Sample/ack
      -- 
    ack_828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_415_index_offset_ack_0, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	514 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (11) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_root_address_calculated
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_offset_calculated
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_Update/ack
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_base_plus_offset/$entry
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_base_plus_offset/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_base_plus_offset/sum_rename_req
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_base_plus_offset/sum_rename_ack
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_request/$entry
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_request/req
      -- 
    ack_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_415_index_offset_ack_1, ack => convTranspose_CP_39_elements(97)); -- 
    req_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(97), ack => addr_of_416_final_reg_req_0); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_request/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_request/ack
      -- 
    ack_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_416_final_reg_ack_0, ack => convTranspose_CP_39_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	514 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	132 
    -- CP-element group 99:  members (19) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_addr_resize/base_resize_ack
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_addr_resize/base_resize_req
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_addr_resize/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_addr_resize/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_address_resized
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_root_address_calculated
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_word_address_calculated
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_address_calculated
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_plus_offset/sum_rename_ack
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_plus_offset/sum_rename_req
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_plus_offset/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_base_plus_offset/$entry
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_word_addrgen/root_register_ack
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_word_addrgen/root_register_req
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_complete/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_complete/ack
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_word_addrgen/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_word_addrgen/$entry
      -- 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_416_final_reg_ack_1, ack => convTranspose_CP_39_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	514 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_update_start_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_Update/cr
      -- 
    ra_857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_419_inst_ack_0, ack => convTranspose_CP_39_elements(100)); -- 
    cr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(100), ack => RPIPE_ConvTranspose_input_pipe_419_inst_req_1); -- 
    -- CP-element group 101:  fork  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (9) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_Sample/rr
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_Sample/rr
      -- 
    ca_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_419_inst_ack_1, ack => convTranspose_CP_39_elements(101)); -- 
    rr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(101), ack => type_cast_423_inst_req_0); -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(101), ack => RPIPE_ConvTranspose_input_pipe_432_inst_req_0); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_Sample/ra
      -- 
    ra_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_423_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	514 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	132 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_Update/ca
      -- 
    ca_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_423_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	101 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_update_start_
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_Update/cr
      -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_432_inst_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    cr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(104), ack => RPIPE_ConvTranspose_input_pipe_432_inst_req_1); -- 
    -- CP-element group 105:  fork  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (9) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_432_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_Sample/rr
      -- 
    ca_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_432_inst_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    rr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(105), ack => type_cast_436_inst_req_0); -- 
    rr_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(105), ack => RPIPE_ConvTranspose_input_pipe_450_inst_req_0); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_Sample/ra
      -- 
    ra_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_436_inst_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	514 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	132 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_Update/ca
      -- 
    ca_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_436_inst_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (6) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_update_start_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_Update/cr
      -- 
    ra_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_450_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    cr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(108), ack => RPIPE_ConvTranspose_input_pipe_450_inst_req_1); -- 
    -- CP-element group 109:  fork  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_450_Update/ca
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_Sample/rr
      -- 
    ca_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_450_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(109), ack => type_cast_454_inst_req_0); -- 
    rr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(109), ack => RPIPE_ConvTranspose_input_pipe_468_inst_req_0); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_Sample/ra
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_454_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	514 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	132 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_Update/ca
      -- 
    ca_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_454_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_update_start_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_Update/cr
      -- 
    ra_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_468_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    cr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(112), ack => RPIPE_ConvTranspose_input_pipe_468_inst_req_1); -- 
    -- CP-element group 113:  fork  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	116 
    -- CP-element group 113:  members (9) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_468_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_Sample/rr
      -- 
    ca_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_468_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    rr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(113), ack => type_cast_472_inst_req_0); -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(113), ack => RPIPE_ConvTranspose_input_pipe_486_inst_req_0); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_Sample/ra
      -- 
    ra_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_472_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	514 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	132 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_update_completed_
      -- 
    ca_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_472_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    -- CP-element group 116:  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	113 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (6) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_update_start_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_sample_completed_
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_486_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(116), ack => RPIPE_ConvTranspose_input_pipe_486_inst_req_1); -- 
    -- CP-element group 117:  fork  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117: 	120 
    -- CP-element group 117:  members (9) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_486_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_sample_start_
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_486_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    rr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(117), ack => type_cast_490_inst_req_0); -- 
    rr_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(117), ack => RPIPE_ConvTranspose_input_pipe_504_inst_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_sample_completed_
      -- 
    ra_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_490_inst_ack_0, ack => convTranspose_CP_39_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	514 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	132 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_Update/$exit
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_490_inst_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	117 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_Update/cr
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_update_start_
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_sample_completed_
      -- 
    ra_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_504_inst_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    cr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(120), ack => RPIPE_ConvTranspose_input_pipe_504_inst_req_1); -- 
    -- CP-element group 121:  fork  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (9) 
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_Update/ca
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_504_update_completed_
      -- 
    ca_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_504_inst_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_508_inst_req_0); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => RPIPE_ConvTranspose_input_pipe_522_inst_req_0); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_sample_completed_
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_508_inst_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	514 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	132 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_update_completed_
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_508_inst_ack_1, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (6) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_Sample/ra
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_update_start_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_sample_completed_
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_522_inst_ack_0, ack => convTranspose_CP_39_elements(124)); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(124), ack => RPIPE_ConvTranspose_input_pipe_522_inst_req_1); -- 
    -- CP-element group 125:  fork  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125: 	128 
    -- CP-element group 125:  members (9) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_Sample/rr
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_Sample/rr
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_522_update_completed_
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_522_inst_ack_1, ack => convTranspose_CP_39_elements(125)); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(125), ack => type_cast_526_inst_req_0); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(125), ack => RPIPE_ConvTranspose_input_pipe_540_inst_req_0); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_Sample/ra
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_Sample/$exit
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_526_inst_ack_0, ack => convTranspose_CP_39_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	514 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	132 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_update_completed_
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_526_inst_ack_1, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	125 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_Update/cr
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_Sample/ra
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_update_start_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_sample_completed_
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_540_inst_ack_0, ack => convTranspose_CP_39_elements(128)); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(128), ack => RPIPE_ConvTranspose_input_pipe_540_inst_req_1); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_Update/ca
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_540_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_Sample/rr
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_Sample/$entry
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_540_inst_ack_1, ack => convTranspose_CP_39_elements(129)); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => type_cast_544_inst_req_0); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_Sample/ra
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_Sample/$exit
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_544_inst_ack_0, ack => convTranspose_CP_39_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	514 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_update_completed_
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_544_inst_ack_1, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	99 
    -- CP-element group 132: 	103 
    -- CP-element group 132: 	107 
    -- CP-element group 132: 	111 
    -- CP-element group 132: 	115 
    -- CP-element group 132: 	119 
    -- CP-element group 132: 	123 
    -- CP-element group 132: 	127 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (9) 
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/word_access_start/word_0/rr
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/word_access_start/word_0/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/word_access_start/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/ptr_deref_552_Split/split_ack
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/ptr_deref_552_Split/split_req
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/ptr_deref_552_Split/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/ptr_deref_552_Split/$entry
      -- 
    rr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(132), ack => ptr_deref_552_store_0_req_0); -- 
    convTranspose_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(99) & convTranspose_CP_39_elements(103) & convTranspose_CP_39_elements(107) & convTranspose_CP_39_elements(111) & convTranspose_CP_39_elements(115) & convTranspose_CP_39_elements(119) & convTranspose_CP_39_elements(123) & convTranspose_CP_39_elements(127) & convTranspose_CP_39_elements(131);
      gj_convTranspose_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/word_access_start/word_0/ra
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/word_access_start/word_0/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/word_access_start/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Sample/$exit
      -- 
    ra_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_552_store_0_ack_0, ack => convTranspose_CP_39_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	514 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (5) 
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Update/word_access_complete/word_0/ca
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Update/word_access_complete/word_0/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Update/word_access_complete/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Update/$exit
      -- 
    ca_1122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_552_store_0_ack_1, ack => convTranspose_CP_39_elements(134)); -- 
    -- CP-element group 135:  branch  join  transition  place  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	96 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (10) 
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565__exit__
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_566__entry__
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_566_dead_link/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_566_else_link/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_566_if_link/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/R_exitcond3_567_place
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_566_eval_test/branch_req
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_566_eval_test/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_566_eval_test/$entry
      -- 
    branch_req_1130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(135), ack => if_stmt_566_branch_req_0); -- 
    convTranspose_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(96) & convTranspose_CP_39_elements(134);
      gj_convTranspose_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  merge  transition  place  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	508 
    -- CP-element group 136:  members (13) 
      -- CP-element group 136: 	 branch_block_stmt_32/merge_stmt_356__exit__
      -- CP-element group 136: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 136: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 136: 	 branch_block_stmt_32/if_stmt_566_if_link/if_choice_transition
      -- CP-element group 136: 	 branch_block_stmt_32/if_stmt_566_if_link/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 136: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/merge_stmt_356_PhiReqMerge
      -- CP-element group 136: 	 branch_block_stmt_32/merge_stmt_356_PhiAck/$entry
      -- CP-element group 136: 	 branch_block_stmt_32/merge_stmt_356_PhiAck/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/merge_stmt_356_PhiAck/dummy
      -- CP-element group 136: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 136: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_566_branch_ack_1, ack => convTranspose_CP_39_elements(136)); -- 
    -- CP-element group 137:  fork  transition  place  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	510 
    -- CP-element group 137: 	511 
    -- CP-element group 137:  members (12) 
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 137: 	 branch_block_stmt_32/if_stmt_566_else_link/else_choice_transition
      -- CP-element group 137: 	 branch_block_stmt_32/if_stmt_566_else_link/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/Sample/rr
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_566_branch_ack_0, ack => convTranspose_CP_39_elements(137)); -- 
    rr_3856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => type_cast_409_inst_req_0); -- 
    cr_3861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => type_cast_409_inst_req_1); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	92 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_sample_completed_
      -- 
    ra_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => convTranspose_CP_39_elements(138)); -- 
    -- CP-element group 139:  transition  place  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	92 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	515 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607__exit__
      -- CP-element group 139: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/type_cast_593_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_578_to_assign_stmt_607/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196_PhiReq/phi_stmt_610/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/$entry
      -- 
    ca_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_1, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	520 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	179 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_Sample/ack
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_sample_complete
      -- 
    ack_1187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_622_index_offset_ack_0, ack => convTranspose_CP_39_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	520 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_request/req
      -- 
    ack_1192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_622_index_offset_ack_1, ack => convTranspose_CP_39_elements(141)); -- 
    req_1201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(141), ack => addr_of_623_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_request/ack
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_request/$exit
      -- 
    ack_1202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_623_final_reg_ack_0, ack => convTranspose_CP_39_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	520 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	176 
    -- CP-element group 143:  members (19) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_word_addrgen/root_register_ack
      -- 
    ack_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_623_final_reg_ack_1, ack => convTranspose_CP_39_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	520 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (6) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_Update/cr
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_Sample/ra
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_update_start_
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_sample_completed_
      -- 
    ra_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_626_inst_ack_0, ack => convTranspose_CP_39_elements(144)); -- 
    cr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(144), ack => RPIPE_ConvTranspose_input_pipe_626_inst_req_1); -- 
    -- CP-element group 145:  fork  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145: 	148 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_Sample/rr
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_Update/ca
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_Sample/rr
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_Sample/$entry
      -- 
    ca_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_626_inst_ack_1, ack => convTranspose_CP_39_elements(145)); -- 
    rr_1229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => type_cast_630_inst_req_0); -- 
    rr_1243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => RPIPE_ConvTranspose_input_pipe_639_inst_req_0); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_Sample/$exit
      -- 
    ra_1230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_630_inst_ack_0, ack => convTranspose_CP_39_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	520 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	176 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_update_completed_
      -- 
    ca_1235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_630_inst_ack_1, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	145 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (6) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_update_start_
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_Update/cr
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_Sample/ra
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_sample_completed_
      -- 
    ra_1244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_639_inst_ack_0, ack => convTranspose_CP_39_elements(148)); -- 
    cr_1248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(148), ack => RPIPE_ConvTranspose_input_pipe_639_inst_req_1); -- 
    -- CP-element group 149:  fork  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149: 	152 
    -- CP-element group 149:  members (9) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_Update/ca
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_639_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_sample_start_
      -- 
    ca_1249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_639_inst_ack_1, ack => convTranspose_CP_39_elements(149)); -- 
    rr_1257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => type_cast_643_inst_req_0); -- 
    rr_1271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => RPIPE_ConvTranspose_input_pipe_657_inst_req_0); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_sample_completed_
      -- 
    ra_1258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_0, ack => convTranspose_CP_39_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	520 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	176 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_update_completed_
      -- 
    ca_1263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_1, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	149 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_Update/cr
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_update_start_
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_sample_completed_
      -- 
    ra_1272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_657_inst_ack_0, ack => convTranspose_CP_39_elements(152)); -- 
    cr_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(152), ack => RPIPE_ConvTranspose_input_pipe_657_inst_req_1); -- 
    -- CP-element group 153:  fork  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	156 
    -- CP-element group 153:  members (9) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_657_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_Sample/rr
      -- 
    ca_1277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_657_inst_ack_1, ack => convTranspose_CP_39_elements(153)); -- 
    rr_1285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => type_cast_661_inst_req_0); -- 
    rr_1299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_675_inst_req_0); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_Sample/ra
      -- 
    ra_1286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_661_inst_ack_0, ack => convTranspose_CP_39_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	520 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	176 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_Update/$exit
      -- 
    ca_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_661_inst_ack_1, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	153 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (6) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_update_start_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_sample_completed_
      -- 
    ra_1300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_675_inst_ack_0, ack => convTranspose_CP_39_elements(156)); -- 
    cr_1304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(156), ack => RPIPE_ConvTranspose_input_pipe_675_inst_req_1); -- 
    -- CP-element group 157:  fork  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: 	160 
    -- CP-element group 157:  members (9) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_Sample/rr
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_675_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_Sample/rr
      -- 
    ca_1305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_675_inst_ack_1, ack => convTranspose_CP_39_elements(157)); -- 
    rr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => type_cast_679_inst_req_0); -- 
    rr_1327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_693_inst_req_0); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_sample_completed_
      -- 
    ra_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_0, ack => convTranspose_CP_39_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	520 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	176 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_update_completed_
      -- 
    ca_1319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_1, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	157 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (6) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_update_start_
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_Sample/ra
      -- 
    ra_1328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_693_inst_ack_0, ack => convTranspose_CP_39_elements(160)); -- 
    cr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(160), ack => RPIPE_ConvTranspose_input_pipe_693_inst_req_1); -- 
    -- CP-element group 161:  fork  transition  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: 	164 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_Sample/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_Sample/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_693_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_Sample/$entry
      -- 
    ca_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_693_inst_ack_1, ack => convTranspose_CP_39_elements(161)); -- 
    rr_1341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => type_cast_697_inst_req_0); -- 
    rr_1355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => RPIPE_ConvTranspose_input_pipe_711_inst_req_0); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_Sample/ra
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_Sample/$exit
      -- 
    ra_1342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_697_inst_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	520 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	176 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_Update/$exit
      -- 
    ca_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_697_inst_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	161 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_Update/cr
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_Sample/ra
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_update_start_
      -- 
    ra_1356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_711_inst_ack_0, ack => convTranspose_CP_39_elements(164)); -- 
    cr_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => RPIPE_ConvTranspose_input_pipe_711_inst_req_1); -- 
    -- CP-element group 165:  fork  transition  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	168 
    -- CP-element group 165:  members (9) 
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_711_update_completed_
      -- 
    ca_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_711_inst_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    rr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(165), ack => type_cast_715_inst_req_0); -- 
    rr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(165), ack => RPIPE_ConvTranspose_input_pipe_729_inst_req_0); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_Sample/$exit
      -- 
    ra_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_715_inst_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	520 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	176 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_Update/$exit
      -- 
    ca_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_715_inst_ack_1, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	165 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_Sample/ra
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_update_start_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_sample_completed_
      -- 
    ra_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_729_inst_ack_0, ack => convTranspose_CP_39_elements(168)); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(168), ack => RPIPE_ConvTranspose_input_pipe_729_inst_req_1); -- 
    -- CP-element group 169:  fork  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	172 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (9) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_Sample/rr
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_729_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_Sample/rr
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_729_inst_ack_1, ack => convTranspose_CP_39_elements(169)); -- 
    rr_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(169), ack => type_cast_733_inst_req_0); -- 
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(169), ack => RPIPE_ConvTranspose_input_pipe_747_inst_req_0); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_sample_completed_
      -- 
    ra_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_733_inst_ack_0, ack => convTranspose_CP_39_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	520 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	176 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_update_completed_
      -- 
    ca_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_733_inst_ack_1, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	169 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_Sample/ra
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_update_start_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_sample_completed_
      -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_747_inst_ack_0, ack => convTranspose_CP_39_elements(172)); -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(172), ack => RPIPE_ConvTranspose_input_pipe_747_inst_req_1); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_747_Update/ca
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_Sample/rr
      -- 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_747_inst_ack_1, ack => convTranspose_CP_39_elements(173)); -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => type_cast_751_inst_req_0); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_Sample/ra
      -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_0, ack => convTranspose_CP_39_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	520 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_Update/ca
      -- 
    ca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_1, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: 	171 
    -- CP-element group 176: 	155 
    -- CP-element group 176: 	159 
    -- CP-element group 176: 	163 
    -- CP-element group 176: 	167 
    -- CP-element group 176: 	151 
    -- CP-element group 176: 	143 
    -- CP-element group 176: 	147 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/ptr_deref_759_Split/$entry
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/ptr_deref_759_Split/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/ptr_deref_759_Split/split_req
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/ptr_deref_759_Split/split_ack
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/word_access_start/$entry
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/word_access_start/word_0/$entry
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/word_access_start/word_0/rr
      -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(176), ack => ptr_deref_759_store_0_req_0); -- 
    convTranspose_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(175) & convTranspose_CP_39_elements(171) & convTranspose_CP_39_elements(155) & convTranspose_CP_39_elements(159) & convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(167) & convTranspose_CP_39_elements(151) & convTranspose_CP_39_elements(143) & convTranspose_CP_39_elements(147);
      gj_convTranspose_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (5) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/word_access_start/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/word_access_start/word_0/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Sample/word_access_start/word_0/ra
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_759_store_0_ack_0, ack => convTranspose_CP_39_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	520 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (5) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Update/word_access_complete/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Update/word_access_complete/word_0/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Update/word_access_complete/word_0/ca
      -- 
    ca_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_759_store_0_ack_1, ack => convTranspose_CP_39_elements(178)); -- 
    -- CP-element group 179:  branch  join  transition  place  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: 	140 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (10) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772__exit__
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_773__entry__
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_773_dead_link/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_773_eval_test/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_773_eval_test/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_773_eval_test/branch_req
      -- CP-element group 179: 	 branch_block_stmt_32/R_exitcond2_774_place
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_773_if_link/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/if_stmt_773_else_link/$entry
      -- 
    branch_req_1489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(179), ack => if_stmt_773_branch_req_0); -- 
    convTranspose_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(178) & convTranspose_CP_39_elements(140);
      gj_convTranspose_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  merge  transition  place  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	521 
    -- CP-element group 180:  members (13) 
      -- CP-element group 180: 	 branch_block_stmt_32/merge_stmt_779__exit__
      -- CP-element group 180: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 180: 	 branch_block_stmt_32/if_stmt_773_if_link/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/if_stmt_773_if_link/if_choice_transition
      -- CP-element group 180: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 180: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 180: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/merge_stmt_779_PhiReqMerge
      -- CP-element group 180: 	 branch_block_stmt_32/merge_stmt_779_PhiAck/$entry
      -- CP-element group 180: 	 branch_block_stmt_32/merge_stmt_779_PhiAck/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/merge_stmt_779_PhiAck/dummy
      -- CP-element group 180: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 180: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_773_branch_ack_1, ack => convTranspose_CP_39_elements(180)); -- 
    -- CP-element group 181:  fork  transition  place  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	516 
    -- CP-element group 181: 	517 
    -- CP-element group 181:  members (12) 
      -- CP-element group 181: 	 branch_block_stmt_32/if_stmt_773_else_link/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/if_stmt_773_else_link/else_choice_transition
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_773_branch_ack_0, ack => convTranspose_CP_39_elements(181)); -- 
    rr_3910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => type_cast_616_inst_req_0); -- 
    cr_3915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => type_cast_616_inst_req_1); -- 
    -- CP-element group 182:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	521 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (18) 
      -- CP-element group 182: 	 branch_block_stmt_32/merge_stmt_804__exit__
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839__entry__
      -- CP-element group 182: 	 branch_block_stmt_32/if_stmt_798_if_link/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/if_stmt_798_if_link/if_choice_transition
      -- CP-element group 182: 	 branch_block_stmt_32/forx_xend250_bbx_xnph757
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_update_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_Update/cr
      -- CP-element group 182: 	 branch_block_stmt_32/forx_xend250_bbx_xnph757_PhiReq/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/forx_xend250_bbx_xnph757_PhiReq/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/merge_stmt_804_PhiReqMerge
      -- CP-element group 182: 	 branch_block_stmt_32/merge_stmt_804_PhiAck/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/merge_stmt_804_PhiAck/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/merge_stmt_804_PhiAck/dummy
      -- 
    if_choice_transition_1516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_798_branch_ack_1, ack => convTranspose_CP_39_elements(182)); -- 
    rr_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_825_inst_req_0); -- 
    cr_1538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(182), ack => type_cast_825_inst_req_1); -- 
    -- CP-element group 183:  transition  place  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	521 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	528 
    -- CP-element group 183:  members (5) 
      -- CP-element group 183: 	 branch_block_stmt_32/if_stmt_798_else_link/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/if_stmt_798_else_link/else_choice_transition
      -- CP-element group 183: 	 branch_block_stmt_32/forx_xend250_forx_xend273
      -- CP-element group 183: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$entry
      -- 
    else_choice_transition_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_798_branch_ack_0, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_Sample/ra
      -- 
    ra_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_825_inst_ack_0, ack => convTranspose_CP_39_elements(184)); -- 
    -- CP-element group 185:  transition  place  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	522 
    -- CP-element group 185:  members (9) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839__exit__
      -- CP-element group 185: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_810_to_assign_stmt_839/type_cast_825_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266_PhiReq/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266_PhiReq/phi_stmt_842/$entry
      -- CP-element group 185: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/$entry
      -- 
    ca_1539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_825_inst_ack_1, ack => convTranspose_CP_39_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	527 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	192 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_sample_complete
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_Sample/ack
      -- 
    ack_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_854_index_offset_ack_0, ack => convTranspose_CP_39_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	527 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (11) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_root_address_calculated
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_offset_calculated
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_Update/ack
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_base_plus_offset/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_base_plus_offset/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_base_plus_offset/sum_rename_req
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_base_plus_offset/sum_rename_ack
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_request/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_request/req
      -- 
    ack_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_854_index_offset_ack_1, ack => convTranspose_CP_39_elements(187)); -- 
    req_1582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(187), ack => addr_of_855_final_reg_req_0); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_request/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_request/ack
      -- 
    ack_1583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_855_final_reg_ack_0, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  join  fork  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	527 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (28) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_complete/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_complete/ack
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_address_calculated
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_word_address_calculated
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_root_address_calculated
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_address_resized
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_addr_resize/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_addr_resize/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_addr_resize/base_resize_req
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_addr_resize/base_resize_ack
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_plus_offset/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_plus_offset/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_plus_offset/sum_rename_req
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_base_plus_offset/sum_rename_ack
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_word_addrgen/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_word_addrgen/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_word_addrgen/root_register_req
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_word_addrgen/root_register_ack
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/ptr_deref_858_Split/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/ptr_deref_858_Split/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/ptr_deref_858_Split/split_req
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/ptr_deref_858_Split/split_ack
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/word_access_start/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/word_access_start/word_0/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/word_access_start/word_0/rr
      -- 
    ack_1588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_855_final_reg_ack_1, ack => convTranspose_CP_39_elements(189)); -- 
    rr_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => ptr_deref_858_store_0_req_0); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (5) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/word_access_start/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/word_access_start/word_0/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Sample/word_access_start/word_0/ra
      -- 
    ra_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_858_store_0_ack_0, ack => convTranspose_CP_39_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	527 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (5) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Update/word_access_complete/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Update/word_access_complete/word_0/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Update/word_access_complete/word_0/ca
      -- 
    ca_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_858_store_0_ack_1, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  branch  join  transition  place  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	186 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (10) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872__exit__
      -- CP-element group 192: 	 branch_block_stmt_32/if_stmt_873__entry__
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/if_stmt_873_dead_link/$entry
      -- CP-element group 192: 	 branch_block_stmt_32/if_stmt_873_eval_test/$entry
      -- CP-element group 192: 	 branch_block_stmt_32/if_stmt_873_eval_test/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/if_stmt_873_eval_test/branch_req
      -- CP-element group 192: 	 branch_block_stmt_32/R_exitcond_874_place
      -- CP-element group 192: 	 branch_block_stmt_32/if_stmt_873_if_link/$entry
      -- CP-element group 192: 	 branch_block_stmt_32/if_stmt_873_else_link/$entry
      -- 
    branch_req_1646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(192), ack => if_stmt_873_branch_req_0); -- 
    convTranspose_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(186) & convTranspose_CP_39_elements(191);
      gj_convTranspose_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  merge  transition  place  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	528 
    -- CP-element group 193:  members (13) 
      -- CP-element group 193: 	 branch_block_stmt_32/merge_stmt_879__exit__
      -- CP-element group 193: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 193: 	 branch_block_stmt_32/if_stmt_873_if_link/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/if_stmt_873_if_link/if_choice_transition
      -- CP-element group 193: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 193: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 193: 	 branch_block_stmt_32/merge_stmt_879_PhiAck/dummy
      -- CP-element group 193: 	 branch_block_stmt_32/merge_stmt_879_PhiAck/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 193: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/merge_stmt_879_PhiReqMerge
      -- CP-element group 193: 	 branch_block_stmt_32/merge_stmt_879_PhiAck/$entry
      -- 
    if_choice_transition_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_873_branch_ack_1, ack => convTranspose_CP_39_elements(193)); -- 
    -- CP-element group 194:  fork  transition  place  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	523 
    -- CP-element group 194: 	524 
    -- CP-element group 194:  members (12) 
      -- CP-element group 194: 	 branch_block_stmt_32/if_stmt_873_else_link/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/if_stmt_873_else_link/else_choice_transition
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_873_branch_ack_0, ack => convTranspose_CP_39_elements(194)); -- 
    rr_3987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_848_inst_req_0); -- 
    cr_3992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(194), ack => type_cast_848_inst_req_1); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	528 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_Sample/cra
      -- 
    cra_1669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_884_call_ack_0, ack => convTranspose_CP_39_elements(195)); -- 
    -- CP-element group 196:  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	528 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (6) 
      -- CP-element group 196: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_Update/cca
      -- CP-element group 196: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_Sample/rr
      -- 
    cca_1674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_884_call_ack_1, ack => convTranspose_CP_39_elements(196)); -- 
    rr_1682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(196), ack => type_cast_889_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_Sample/ra
      -- 
    ra_1683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_889_inst_ack_0, ack => convTranspose_CP_39_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	528 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	449 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_Update/ca
      -- 
    ca_1688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_889_inst_ack_1, ack => convTranspose_CP_39_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	528 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_update_start_
      -- CP-element group 199: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_Sample/ack
      -- CP-element group 199: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_Update/req
      -- 
    ack_1697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_891_inst_ack_0, ack => convTranspose_CP_39_elements(199)); -- 
    req_1701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(199), ack => WPIPE_Block0_start_891_inst_req_1); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_Update/ack
      -- CP-element group 200: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_Sample/req
      -- 
    ack_1702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_891_inst_ack_1, ack => convTranspose_CP_39_elements(200)); -- 
    req_1710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(200), ack => WPIPE_Block0_start_894_inst_req_0); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_update_start_
      -- CP-element group 201: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_Update/req
      -- 
    ack_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_894_inst_ack_0, ack => convTranspose_CP_39_elements(201)); -- 
    req_1715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(201), ack => WPIPE_Block0_start_894_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_894_Update/ack
      -- CP-element group 202: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_Sample/req
      -- 
    ack_1716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_894_inst_ack_1, ack => convTranspose_CP_39_elements(202)); -- 
    req_1724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => WPIPE_Block0_start_897_inst_req_0); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_update_start_
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_Sample/ack
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_Update/req
      -- 
    ack_1725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_897_inst_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    req_1729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(203), ack => WPIPE_Block0_start_897_inst_req_1); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_897_Update/ack
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_Sample/req
      -- 
    ack_1730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_897_inst_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    req_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(204), ack => WPIPE_Block0_start_900_inst_req_0); -- 
    -- CP-element group 205:  transition  input  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (6) 
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_update_start_
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_Sample/ack
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_Update/$entry
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_Update/req
      -- 
    ack_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_900_inst_ack_0, ack => convTranspose_CP_39_elements(205)); -- 
    req_1743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(205), ack => WPIPE_Block0_start_900_inst_req_1); -- 
    -- CP-element group 206:  transition  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (6) 
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_900_Update/ack
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_Sample/req
      -- 
    ack_1744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_900_inst_ack_1, ack => convTranspose_CP_39_elements(206)); -- 
    req_1752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(206), ack => WPIPE_Block0_start_903_inst_req_0); -- 
    -- CP-element group 207:  transition  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (6) 
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_update_start_
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_Sample/ack
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_Update/req
      -- 
    ack_1753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_903_inst_ack_0, ack => convTranspose_CP_39_elements(207)); -- 
    req_1757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(207), ack => WPIPE_Block0_start_903_inst_req_1); -- 
    -- CP-element group 208:  transition  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_903_Update/ack
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_Sample/req
      -- 
    ack_1758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_903_inst_ack_1, ack => convTranspose_CP_39_elements(208)); -- 
    req_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => WPIPE_Block0_start_906_inst_req_0); -- 
    -- CP-element group 209:  transition  input  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (6) 
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_update_start_
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_Sample/ack
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_Update/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_Update/req
      -- 
    ack_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_906_inst_ack_0, ack => convTranspose_CP_39_elements(209)); -- 
    req_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(209), ack => WPIPE_Block0_start_906_inst_req_1); -- 
    -- CP-element group 210:  transition  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (6) 
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_906_Update/ack
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_Sample/req
      -- 
    ack_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_906_inst_ack_1, ack => convTranspose_CP_39_elements(210)); -- 
    req_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => WPIPE_Block0_start_909_inst_req_0); -- 
    -- CP-element group 211:  transition  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211:  members (6) 
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_update_start_
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_Sample/ack
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_Update/req
      -- 
    ack_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_909_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    req_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(211), ack => WPIPE_Block0_start_909_inst_req_1); -- 
    -- CP-element group 212:  transition  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (6) 
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_909_Update/ack
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_Sample/req
      -- 
    ack_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_909_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    req_1794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(212), ack => WPIPE_Block0_start_912_inst_req_0); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_update_start_
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_Sample/ack
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_Update/req
      -- 
    ack_1795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_912_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    req_1799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(213), ack => WPIPE_Block0_start_912_inst_req_1); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_912_Update/ack
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_Sample/req
      -- 
    ack_1800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_912_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    req_1808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(214), ack => WPIPE_Block0_start_915_inst_req_0); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_update_start_
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_Update/req
      -- 
    ack_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_915_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    req_1813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(215), ack => WPIPE_Block0_start_915_inst_req_1); -- 
    -- CP-element group 216:  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_915_Update/ack
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_Sample/req
      -- 
    ack_1814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_915_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    req_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(216), ack => WPIPE_Block0_start_918_inst_req_0); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_update_start_
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_Sample/ack
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_Update/req
      -- 
    ack_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_918_inst_ack_0, ack => convTranspose_CP_39_elements(217)); -- 
    req_1827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => WPIPE_Block0_start_918_inst_req_1); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (6) 
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_918_Update/ack
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_Sample/req
      -- 
    ack_1828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_918_inst_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    req_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => WPIPE_Block0_start_921_inst_req_0); -- 
    -- CP-element group 219:  transition  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (6) 
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_update_start_
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_Sample/ack
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_Update/req
      -- 
    ack_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_921_inst_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(219), ack => WPIPE_Block0_start_921_inst_req_1); -- 
    -- CP-element group 220:  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (6) 
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_921_Update/ack
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_Sample/req
      -- 
    ack_1842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_921_inst_ack_1, ack => convTranspose_CP_39_elements(220)); -- 
    req_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(220), ack => WPIPE_Block0_start_924_inst_req_0); -- 
    -- CP-element group 221:  transition  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (6) 
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_update_start_
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_Sample/ack
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_Update/req
      -- 
    ack_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_924_inst_ack_0, ack => convTranspose_CP_39_elements(221)); -- 
    req_1855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(221), ack => WPIPE_Block0_start_924_inst_req_1); -- 
    -- CP-element group 222:  transition  input  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (6) 
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_924_Update/ack
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_Sample/req
      -- 
    ack_1856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_924_inst_ack_1, ack => convTranspose_CP_39_elements(222)); -- 
    req_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(222), ack => WPIPE_Block0_start_927_inst_req_0); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (6) 
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_update_start_
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_Update/req
      -- 
    ack_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_927_inst_ack_0, ack => convTranspose_CP_39_elements(223)); -- 
    req_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => WPIPE_Block0_start_927_inst_req_1); -- 
    -- CP-element group 224:  transition  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (6) 
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_927_Update/ack
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_sample_start_
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_Sample/req
      -- 
    ack_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_927_inst_ack_1, ack => convTranspose_CP_39_elements(224)); -- 
    req_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(224), ack => WPIPE_Block0_start_930_inst_req_0); -- 
    -- CP-element group 225:  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (6) 
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_update_start_
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_Sample/ack
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_Update/req
      -- 
    ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_930_inst_ack_0, ack => convTranspose_CP_39_elements(225)); -- 
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => WPIPE_Block0_start_930_inst_req_1); -- 
    -- CP-element group 226:  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (6) 
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_930_Update/ack
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_Sample/req
      -- 
    ack_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_930_inst_ack_1, ack => convTranspose_CP_39_elements(226)); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(226), ack => WPIPE_Block0_start_933_inst_req_0); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (6) 
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_update_start_
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_Sample/ack
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_Update/req
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_933_inst_ack_0, ack => convTranspose_CP_39_elements(227)); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(227), ack => WPIPE_Block0_start_933_inst_req_1); -- 
    -- CP-element group 228:  transition  input  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (6) 
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_933_Update/ack
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_Sample/req
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_933_inst_ack_1, ack => convTranspose_CP_39_elements(228)); -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => WPIPE_Block0_start_936_inst_req_0); -- 
    -- CP-element group 229:  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (6) 
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_sample_completed_
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_update_start_
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_Sample/ack
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_Update/req
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_936_inst_ack_0, ack => convTranspose_CP_39_elements(229)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(229), ack => WPIPE_Block0_start_936_inst_req_1); -- 
    -- CP-element group 230:  transition  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (6) 
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_936_Update/ack
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_Sample/req
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_936_inst_ack_1, ack => convTranspose_CP_39_elements(230)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => WPIPE_Block0_start_939_inst_req_0); -- 
    -- CP-element group 231:  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (6) 
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_update_start_
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_Sample/ack
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_Update/req
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_939_inst_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(231), ack => WPIPE_Block0_start_939_inst_req_1); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_939_Update/ack
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_Sample/req
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_939_inst_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(232), ack => WPIPE_Block0_start_942_inst_req_0); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_update_start_
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_Sample/ack
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_Update/req
      -- 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_942_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(233), ack => WPIPE_Block0_start_942_inst_req_1); -- 
    -- CP-element group 234:  transition  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_942_Update/ack
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_Sample/req
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_942_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block0_start_945_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_update_start_
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_Update/req
      -- 
    ack_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_945_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block0_start_945_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_945_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_sample_start_
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_945_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block0_start_949_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_Update/req
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_update_start_
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_949_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block0_start_949_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_949_update_completed_
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_949_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block0_start_953_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_update_start_
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_Update/req
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_Sample/$exit
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block0_start_953_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_Sample/req
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_953_Update/$exit
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block0_start_957_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_Update/req
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_sample_completed_
      -- 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_957_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block0_start_957_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_957_update_completed_
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_957_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block0_start_961_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_update_start_
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_Update/req
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_961_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block0_start_961_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_961_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_Sample/$entry
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_961_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block0_start_964_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_Update/req
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_update_start_
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_sample_completed_
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_964_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block0_start_964_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_964_update_completed_
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_964_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block0_start_967_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_Update/req
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_sample_completed_
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_967_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block0_start_967_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_967_update_completed_
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_967_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block0_start_970_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_Update/req
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_sample_completed_
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_970_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block0_start_970_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_970_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_Sample/req
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_Sample/$entry
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_970_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block0_start_973_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_Update/req
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_update_start_
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_973_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block0_start_973_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_973_update_completed_
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_973_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block0_start_976_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_update_start_
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_Update/req
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_Update/$entry
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block0_start_976_inst_req_1); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	449 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_976_Update/$exit
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_976_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	528 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_Update/req
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_sample_completed_
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_979_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block1_start_979_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_update_completed_
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_979_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block1_start_982_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_Update/req
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_update_start_
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_sample_completed_
      -- 
    ack_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_982_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block1_start_982_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_982_update_completed_
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_982_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    req_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(258), ack => WPIPE_Block1_start_985_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_Update/req
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_sample_completed_
      -- 
    ack_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_985_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block1_start_985_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_985_update_completed_
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_985_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block1_start_988_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_Update/req
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_update_start_
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_sample_completed_
      -- 
    ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_988_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block1_start_988_inst_req_1); -- 
    -- CP-element group 262:  transition  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (6) 
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_Sample/req
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_988_update_completed_
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_988_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    req_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(262), ack => WPIPE_Block1_start_991_inst_req_0); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_update_start_
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_Update/req
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_Sample/ack
      -- 
    ack_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_991_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block1_start_991_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_Sample/req
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_991_update_completed_
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_991_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block1_start_994_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_update_start_
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_Update/req
      -- 
    ack_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_994_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block1_start_994_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_994_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_Sample/req
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_994_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block1_start_997_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_update_start_
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_Update/req
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_Sample/ack
      -- 
    ack_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_997_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block1_start_997_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_997_Update/$exit
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_997_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block1_start_1000_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_Update/req
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_update_start_
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_sample_completed_
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1000_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block1_start_1000_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1000_update_completed_
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1000_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block1_start_1003_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_Update/req
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_update_start_
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_sample_completed_
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1003_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block1_start_1003_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1003_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_Sample/$entry
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1003_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block1_start_1006_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_Update/req
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_update_start_
      -- 
    ack_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1006_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block1_start_1006_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1006_update_completed_
      -- 
    ack_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1006_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block1_start_1009_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_Update/req
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_sample_completed_
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1009_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block1_start_1009_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1009_update_completed_
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1009_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block1_start_1012_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_Update/req
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_update_start_
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_sample_completed_
      -- 
    ack_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1012_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block1_start_1012_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1012_update_completed_
      -- 
    ack_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1012_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block1_start_1015_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_Update/req
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_update_start_
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_Update/$entry
      -- 
    ack_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1015_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block1_start_1015_inst_req_1); -- 
    -- CP-element group 280:  transition  input  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (6) 
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_Sample/req
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1015_Update/ack
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1015_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(280), ack => WPIPE_Block1_start_1018_inst_req_0); -- 
    -- CP-element group 281:  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_Update/req
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_Sample/ack
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_sample_completed_
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1018_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(281), ack => WPIPE_Block1_start_1018_inst_req_1); -- 
    -- CP-element group 282:  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (6) 
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_Update/ack
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_Sample/req
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1018_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_Sample/$entry
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1018_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    req_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(282), ack => WPIPE_Block1_start_1021_inst_req_0); -- 
    -- CP-element group 283:  transition  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (6) 
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_sample_completed_
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_Update/req
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_Sample/ack
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_update_start_
      -- 
    ack_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1021_inst_ack_0, ack => convTranspose_CP_39_elements(283)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block1_start_1021_inst_req_1); -- 
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_Update/ack
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_Sample/req
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1021_update_completed_
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1021_inst_ack_1, ack => convTranspose_CP_39_elements(284)); -- 
    req_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(284), ack => WPIPE_Block1_start_1024_inst_req_0); -- 
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_Update/req
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_update_start_
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_Sample/ack
      -- 
    ack_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1024_inst_ack_0, ack => convTranspose_CP_39_elements(285)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(285), ack => WPIPE_Block1_start_1024_inst_req_1); -- 
    -- CP-element group 286:  transition  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (6) 
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1024_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_Sample/req
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_sample_start_
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1024_inst_ack_1, ack => convTranspose_CP_39_elements(286)); -- 
    req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(286), ack => WPIPE_Block1_start_1027_inst_req_0); -- 
    -- CP-element group 287:  transition  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (6) 
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_Update/req
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_Sample/ack
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_sample_completed_
      -- 
    ack_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1027_inst_ack_0, ack => convTranspose_CP_39_elements(287)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(287), ack => WPIPE_Block1_start_1027_inst_req_1); -- 
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_Update/ack
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1027_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_sample_start_
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1027_inst_ack_1, ack => convTranspose_CP_39_elements(288)); -- 
    req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block1_start_1030_inst_req_0); -- 
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_Update/req
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_sample_completed_
      -- 
    ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1030_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block1_start_1030_inst_req_1); -- 
    -- CP-element group 290:  transition  input  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	293 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1030_update_completed_
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1030_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	528 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_Sample/ra
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_sample_completed_
      -- 
    ra_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	528 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_Update/ca
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_update_completed_
      -- 
    ca_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	290 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_sample_start_
      -- 
    req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block1_start_1037_inst_req_0); -- 
    convTranspose_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(290) & convTranspose_CP_39_elements(292);
      gj_convTranspose_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_Update/req
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_Sample/ack
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_update_start_
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_sample_completed_
      -- 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_0, ack => convTranspose_CP_39_elements(294)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block1_start_1037_inst_req_1); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	298 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_Update/ack
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1037_update_completed_
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_1, ack => convTranspose_CP_39_elements(295)); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	528 
    -- CP-element group 296: successors 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_Sample/ra
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_sample_completed_
      -- 
    ra_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1048_inst_ack_0, ack => convTranspose_CP_39_elements(296)); -- 
    -- CP-element group 297:  fork  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	528 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297: 	301 
    -- CP-element group 297: 	304 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_Update/ca
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_update_completed_
      -- 
    ca_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1048_inst_ack_1, ack => convTranspose_CP_39_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	295 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_sample_start_
      -- 
    req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block1_start_1050_inst_req_0); -- 
    convTranspose_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(295) & convTranspose_CP_39_elements(297);
      gj_convTranspose_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_update_start_
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_Update/req
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_Update/$entry
      -- 
    ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1050_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block1_start_1050_inst_req_1); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1050_Update/$exit
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1050_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	297 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_Sample/req
      -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block1_start_1053_inst_req_0); -- 
    convTranspose_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(297) & convTranspose_CP_39_elements(300);
      gj_convTranspose_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_sample_completed_
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_update_start_
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_Sample/$exit
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_Sample/ack
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_Update/req
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_Update/$entry
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1053_inst_ack_0, ack => convTranspose_CP_39_elements(302)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block1_start_1053_inst_req_1); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_update_completed_
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_Update/ack
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1053_Update/$exit
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1053_inst_ack_1, ack => convTranspose_CP_39_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	297 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_Sample/$entry
      -- 
    req_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block1_start_1056_inst_req_0); -- 
    convTranspose_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(297) & convTranspose_CP_39_elements(303);
      gj_convTranspose_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_Update/req
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_update_start_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_Sample/$exit
      -- 
    ack_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1056_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block1_start_1056_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1056_update_completed_
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1056_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(306), ack => WPIPE_Block1_start_1059_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_update_start_
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_Update/req
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1059_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block1_start_1059_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1059_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_Sample/req
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1059_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block1_start_1062_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_update_start_
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_Update/req
      -- 
    ack_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1062_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block1_start_1062_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1062_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_Sample/req
      -- 
    ack_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1062_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(310), ack => WPIPE_Block1_start_1065_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_update_start_
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1065_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => WPIPE_Block1_start_1065_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1065_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_Sample/req
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1065_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    req_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(312), ack => WPIPE_Block1_start_1068_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_update_start_
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_Update/req
      -- 
    ack_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1068_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    req_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => WPIPE_Block1_start_1068_inst_req_1); -- 
    -- CP-element group 314:  transition  input  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (6) 
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1068_Update/ack
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_sample_start_
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_Sample/$entry
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_Sample/req
      -- 
    ack_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1068_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(314), ack => WPIPE_Block1_start_1071_inst_req_0); -- 
    -- CP-element group 315:  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (6) 
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_update_start_
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_Sample/ack
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_Update/req
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1071_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(315), ack => WPIPE_Block1_start_1071_inst_req_1); -- 
    -- CP-element group 316:  transition  input  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (6) 
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1071_Update/ack
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_sample_start_
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_Sample/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1071_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    req_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(316), ack => WPIPE_Block1_start_1074_inst_req_0); -- 
    -- CP-element group 317:  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_sample_completed_
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_update_start_
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_Sample/ack
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_Update/req
      -- 
    ack_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1074_inst_ack_0, ack => convTranspose_CP_39_elements(317)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => WPIPE_Block1_start_1074_inst_req_1); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	449 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_update_completed_
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_1074_Update/ack
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1074_inst_ack_1, ack => convTranspose_CP_39_elements(318)); -- 
    -- CP-element group 319:  transition  input  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	528 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (6) 
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_update_start_
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_Sample/ack
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1077_inst_ack_0, ack => convTranspose_CP_39_elements(319)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(319), ack => WPIPE_Block2_start_1077_inst_req_1); -- 
    -- CP-element group 320:  transition  input  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (6) 
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_Update/ack
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_sample_start_
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_Sample/$entry
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_Sample/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1077_inst_ack_1, ack => convTranspose_CP_39_elements(320)); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(320), ack => WPIPE_Block2_start_1080_inst_req_0); -- 
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_sample_completed_
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_update_start_
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_Sample/ack
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_Update/req
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1080_inst_ack_0, ack => convTranspose_CP_39_elements(321)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(321), ack => WPIPE_Block2_start_1080_inst_req_1); -- 
    -- CP-element group 322:  transition  input  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (6) 
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_update_completed_
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1080_Update/ack
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_Sample/req
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1080_inst_ack_1, ack => convTranspose_CP_39_elements(322)); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(322), ack => WPIPE_Block2_start_1083_inst_req_0); -- 
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_update_start_
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_Update/req
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1083_inst_ack_0, ack => convTranspose_CP_39_elements(323)); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_Block2_start_1083_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1083_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_Sample/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1083_inst_ack_1, ack => convTranspose_CP_39_elements(324)); -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_Block2_start_1086_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_update_start_
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_Update/req
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1086_inst_ack_0, ack => convTranspose_CP_39_elements(325)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => WPIPE_Block2_start_1086_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1086_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_Sample/req
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1086_inst_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => WPIPE_Block2_start_1089_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_update_start_
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_Update/req
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1089_inst_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(327), ack => WPIPE_Block2_start_1089_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1089_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_Sample/req
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1089_inst_ack_1, ack => convTranspose_CP_39_elements(328)); -- 
    req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(328), ack => WPIPE_Block2_start_1092_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_update_start_
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_Update/req
      -- 
    ack_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1092_inst_ack_0, ack => convTranspose_CP_39_elements(329)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(329), ack => WPIPE_Block2_start_1092_inst_req_1); -- 
    -- CP-element group 330:  transition  input  output  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (6) 
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1092_Update/ack
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_sample_start_
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_Sample/$entry
      -- CP-element group 330: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_Sample/req
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1092_inst_ack_1, ack => convTranspose_CP_39_elements(330)); -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(330), ack => WPIPE_Block2_start_1095_inst_req_0); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_update_start_
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_Update/req
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1095_inst_ack_0, ack => convTranspose_CP_39_elements(331)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => WPIPE_Block2_start_1095_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1095_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_Sample/req
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1095_inst_ack_1, ack => convTranspose_CP_39_elements(332)); -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(332), ack => WPIPE_Block2_start_1098_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_update_start_
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_Update/req
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1098_inst_ack_0, ack => convTranspose_CP_39_elements(333)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => WPIPE_Block2_start_1098_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1098_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_Sample/req
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1098_inst_ack_1, ack => convTranspose_CP_39_elements(334)); -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(334), ack => WPIPE_Block2_start_1101_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_update_start_
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_Update/req
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1101_inst_ack_0, ack => convTranspose_CP_39_elements(335)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => WPIPE_Block2_start_1101_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1101_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_Sample/req
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1101_inst_ack_1, ack => convTranspose_CP_39_elements(336)); -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(336), ack => WPIPE_Block2_start_1104_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_update_start_
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_Update/req
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1104_inst_ack_0, ack => convTranspose_CP_39_elements(337)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(337), ack => WPIPE_Block2_start_1104_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1104_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_Sample/req
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1104_inst_ack_1, ack => convTranspose_CP_39_elements(338)); -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(338), ack => WPIPE_Block2_start_1107_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_update_start_
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_Update/req
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1107_inst_ack_0, ack => convTranspose_CP_39_elements(339)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(339), ack => WPIPE_Block2_start_1107_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1107_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_Sample/req
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1107_inst_ack_1, ack => convTranspose_CP_39_elements(340)); -- 
    req_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(340), ack => WPIPE_Block2_start_1110_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_update_start_
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_Update/req
      -- 
    ack_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1110_inst_ack_0, ack => convTranspose_CP_39_elements(341)); -- 
    req_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(341), ack => WPIPE_Block2_start_1110_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1110_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_Sample/req
      -- 
    ack_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1110_inst_ack_1, ack => convTranspose_CP_39_elements(342)); -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(342), ack => WPIPE_Block2_start_1113_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_update_start_
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_Update/req
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_0, ack => convTranspose_CP_39_elements(343)); -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(343), ack => WPIPE_Block2_start_1113_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1113_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_Sample/req
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1113_inst_ack_1, ack => convTranspose_CP_39_elements(344)); -- 
    req_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(344), ack => WPIPE_Block2_start_1116_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_update_start_
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_Update/req
      -- 
    ack_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1116_inst_ack_0, ack => convTranspose_CP_39_elements(345)); -- 
    req_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(345), ack => WPIPE_Block2_start_1116_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1116_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_Sample/req
      -- 
    ack_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1116_inst_ack_1, ack => convTranspose_CP_39_elements(346)); -- 
    req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(346), ack => WPIPE_Block2_start_1119_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_update_start_
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_Update/req
      -- 
    ack_2705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_0, ack => convTranspose_CP_39_elements(347)); -- 
    req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(347), ack => WPIPE_Block2_start_1119_inst_req_1); -- 
    -- CP-element group 348:  transition  input  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (6) 
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1119_Update/ack
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_sample_start_
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_Sample/$entry
      -- CP-element group 348: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_Sample/req
      -- 
    ack_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_1, ack => convTranspose_CP_39_elements(348)); -- 
    req_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(348), ack => WPIPE_Block2_start_1122_inst_req_0); -- 
    -- CP-element group 349:  transition  input  output  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (6) 
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_update_start_
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_Sample/ack
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_Update/$entry
      -- CP-element group 349: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_Update/req
      -- 
    ack_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_0, ack => convTranspose_CP_39_elements(349)); -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(349), ack => WPIPE_Block2_start_1122_inst_req_1); -- 
    -- CP-element group 350:  transition  input  output  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (6) 
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1122_Update/ack
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_sample_start_
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_Sample/req
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_1, ack => convTranspose_CP_39_elements(350)); -- 
    req_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(350), ack => WPIPE_Block2_start_1125_inst_req_0); -- 
    -- CP-element group 351:  transition  input  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (6) 
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_sample_completed_
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_update_start_
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_Sample/ack
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_Update/$entry
      -- CP-element group 351: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_Update/req
      -- 
    ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1125_inst_ack_0, ack => convTranspose_CP_39_elements(351)); -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => WPIPE_Block2_start_1125_inst_req_1); -- 
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_update_completed_
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1125_Update/ack
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_sample_start_
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_Sample/$entry
      -- CP-element group 352: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_Sample/req
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1125_inst_ack_1, ack => convTranspose_CP_39_elements(352)); -- 
    req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_Block2_start_1128_inst_req_0); -- 
    -- CP-element group 353:  transition  input  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (6) 
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_sample_completed_
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_update_start_
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_Sample/$exit
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_Sample/ack
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_Update/req
      -- 
    ack_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1128_inst_ack_0, ack => convTranspose_CP_39_elements(353)); -- 
    req_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(353), ack => WPIPE_Block2_start_1128_inst_req_1); -- 
    -- CP-element group 354:  transition  input  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (6) 
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_update_completed_
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_Update/$exit
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1128_Update/ack
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_Sample/req
      -- 
    ack_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1128_inst_ack_1, ack => convTranspose_CP_39_elements(354)); -- 
    req_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(354), ack => WPIPE_Block2_start_1131_inst_req_0); -- 
    -- CP-element group 355:  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (6) 
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_update_start_
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_Sample/ack
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_Update/req
      -- 
    ack_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1131_inst_ack_0, ack => convTranspose_CP_39_elements(355)); -- 
    req_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => WPIPE_Block2_start_1131_inst_req_1); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	359 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1131_Update/ack
      -- 
    ack_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1131_inst_ack_1, ack => convTranspose_CP_39_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	528 
    -- CP-element group 357: successors 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_Sample/ra
      -- 
    ra_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1143_inst_ack_0, ack => convTranspose_CP_39_elements(357)); -- 
    -- CP-element group 358:  fork  transition  input  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	528 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358: 	362 
    -- CP-element group 358: 	365 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_Update/ca
      -- 
    ca_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1143_inst_ack_1, ack => convTranspose_CP_39_elements(358)); -- 
    -- CP-element group 359:  join  transition  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	356 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_sample_start_
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_Sample/req
      -- 
    req_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(359), ack => WPIPE_Block2_start_1145_inst_req_0); -- 
    convTranspose_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(356) & convTranspose_CP_39_elements(358);
      gj_convTranspose_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_update_start_
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_Sample/ack
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_Update/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_Update/req
      -- 
    ack_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1145_inst_ack_0, ack => convTranspose_CP_39_elements(360)); -- 
    req_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => WPIPE_Block2_start_1145_inst_req_1); -- 
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1145_Update/ack
      -- 
    ack_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1145_inst_ack_1, ack => convTranspose_CP_39_elements(361)); -- 
    -- CP-element group 362:  join  transition  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	358 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_Sample/req
      -- 
    req_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(362), ack => WPIPE_Block2_start_1148_inst_req_0); -- 
    convTranspose_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(358) & convTranspose_CP_39_elements(361);
      gj_convTranspose_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_update_start_
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_Update/req
      -- 
    ack_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1148_inst_ack_0, ack => convTranspose_CP_39_elements(363)); -- 
    req_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(363), ack => WPIPE_Block2_start_1148_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1148_Update/ack
      -- 
    ack_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1148_inst_ack_1, ack => convTranspose_CP_39_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	358 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_Sample/req
      -- 
    req_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(365), ack => WPIPE_Block2_start_1151_inst_req_0); -- 
    convTranspose_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(358) & convTranspose_CP_39_elements(364);
      gj_convTranspose_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  transition  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (6) 
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_sample_completed_
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_update_start_
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_Sample/$exit
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_Sample/ack
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_Update/req
      -- 
    ack_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1151_inst_ack_0, ack => convTranspose_CP_39_elements(366)); -- 
    req_2821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => WPIPE_Block2_start_1151_inst_req_1); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_update_completed_
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_Update/$exit
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1151_Update/ack
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_sample_start_
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_Sample/req
      -- 
    ack_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1151_inst_ack_1, ack => convTranspose_CP_39_elements(367)); -- 
    req_2830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => WPIPE_Block2_start_1154_inst_req_0); -- 
    -- CP-element group 368:  transition  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_update_start_
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_Sample/ack
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_Update/req
      -- 
    ack_2831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1154_inst_ack_0, ack => convTranspose_CP_39_elements(368)); -- 
    req_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(368), ack => WPIPE_Block2_start_1154_inst_req_1); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1154_Update/ack
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_sample_start_
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_Sample/req
      -- 
    ack_2836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1154_inst_ack_1, ack => convTranspose_CP_39_elements(369)); -- 
    req_2844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(369), ack => WPIPE_Block2_start_1157_inst_req_0); -- 
    -- CP-element group 370:  transition  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_update_start_
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_Sample/ack
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_Update/req
      -- 
    ack_2845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1157_inst_ack_0, ack => convTranspose_CP_39_elements(370)); -- 
    req_2849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(370), ack => WPIPE_Block2_start_1157_inst_req_1); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_Sample/req
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1157_Update/ack
      -- CP-element group 371: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_sample_start_
      -- 
    ack_2850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1157_inst_ack_1, ack => convTranspose_CP_39_elements(371)); -- 
    req_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(371), ack => WPIPE_Block2_start_1160_inst_req_0); -- 
    -- CP-element group 372:  transition  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_update_start_
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_Sample/ack
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_Update/req
      -- 
    ack_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1160_inst_ack_0, ack => convTranspose_CP_39_elements(372)); -- 
    req_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => WPIPE_Block2_start_1160_inst_req_1); -- 
    -- CP-element group 373:  transition  input  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (6) 
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1160_Update/ack
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_Sample/req
      -- 
    ack_2864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1160_inst_ack_1, ack => convTranspose_CP_39_elements(373)); -- 
    req_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => WPIPE_Block2_start_1163_inst_req_0); -- 
    -- CP-element group 374:  transition  input  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (6) 
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_update_start_
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_Sample/ack
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_Update/req
      -- 
    ack_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1163_inst_ack_0, ack => convTranspose_CP_39_elements(374)); -- 
    req_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(374), ack => WPIPE_Block2_start_1163_inst_req_1); -- 
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1163_Update/ack
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_Sample/req
      -- 
    ack_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1163_inst_ack_1, ack => convTranspose_CP_39_elements(375)); -- 
    req_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => WPIPE_Block2_start_1166_inst_req_0); -- 
    -- CP-element group 376:  transition  input  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_update_start_
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_Sample/ack
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_Update/req
      -- 
    ack_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1166_inst_ack_0, ack => convTranspose_CP_39_elements(376)); -- 
    req_2891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(376), ack => WPIPE_Block2_start_1166_inst_req_1); -- 
    -- CP-element group 377:  transition  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377:  members (6) 
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1166_Update/ack
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_Sample/req
      -- 
    ack_2892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1166_inst_ack_1, ack => convTranspose_CP_39_elements(377)); -- 
    req_2900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => WPIPE_Block2_start_1169_inst_req_0); -- 
    -- CP-element group 378:  transition  input  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378:  members (6) 
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_update_start_
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_Sample/ack
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_Update/req
      -- 
    ack_2901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1169_inst_ack_0, ack => convTranspose_CP_39_elements(378)); -- 
    req_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(378), ack => WPIPE_Block2_start_1169_inst_req_1); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	378 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	449 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1169_Update/ack
      -- 
    ack_2906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1169_inst_ack_1, ack => convTranspose_CP_39_elements(379)); -- 
    -- CP-element group 380:  transition  input  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	528 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (6) 
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_update_start_
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_Sample/ack
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_Update/req
      -- 
    ack_2915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1172_inst_ack_0, ack => convTranspose_CP_39_elements(380)); -- 
    req_2919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(380), ack => WPIPE_Block3_start_1172_inst_req_1); -- 
    -- CP-element group 381:  transition  input  output  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (6) 
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_Update/ack
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_sample_start_
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_Sample/$entry
      -- CP-element group 381: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_Sample/req
      -- 
    ack_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1172_inst_ack_1, ack => convTranspose_CP_39_elements(381)); -- 
    req_2928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(381), ack => WPIPE_Block3_start_1175_inst_req_0); -- 
    -- CP-element group 382:  transition  input  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (6) 
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_update_start_
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_Sample/ack
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_Update/req
      -- 
    ack_2929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_0, ack => convTranspose_CP_39_elements(382)); -- 
    req_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(382), ack => WPIPE_Block3_start_1175_inst_req_1); -- 
    -- CP-element group 383:  transition  input  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (6) 
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1175_Update/ack
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_Sample/req
      -- 
    ack_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_1, ack => convTranspose_CP_39_elements(383)); -- 
    req_2942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(383), ack => WPIPE_Block3_start_1178_inst_req_0); -- 
    -- CP-element group 384:  transition  input  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (6) 
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_Sample/ack
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_Update/req
      -- 
    ack_2943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    req_2947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => WPIPE_Block3_start_1178_inst_req_1); -- 
    -- CP-element group 385:  transition  input  output  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385:  members (6) 
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1178_Update/ack
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_Sample/req
      -- 
    ack_2948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_1, ack => convTranspose_CP_39_elements(385)); -- 
    req_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(385), ack => WPIPE_Block3_start_1181_inst_req_0); -- 
    -- CP-element group 386:  transition  input  output  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	387 
    -- CP-element group 386:  members (6) 
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_update_start_
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_Sample/ack
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_Update/req
      -- 
    ack_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    req_2961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(386), ack => WPIPE_Block3_start_1181_inst_req_1); -- 
    -- CP-element group 387:  transition  input  output  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	386 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (6) 
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1181_Update/ack
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_sample_start_
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_Sample/$entry
      -- CP-element group 387: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_Sample/req
      -- 
    ack_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_1, ack => convTranspose_CP_39_elements(387)); -- 
    req_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(387), ack => WPIPE_Block3_start_1184_inst_req_0); -- 
    -- CP-element group 388:  transition  input  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (6) 
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_sample_completed_
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_update_start_
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_Sample/ack
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_Update/$entry
      -- CP-element group 388: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_Update/req
      -- 
    ack_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_0, ack => convTranspose_CP_39_elements(388)); -- 
    req_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(388), ack => WPIPE_Block3_start_1184_inst_req_1); -- 
    -- CP-element group 389:  transition  input  output  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (6) 
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_Sample/req
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1184_Update/ack
      -- CP-element group 389: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_sample_start_
      -- 
    ack_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_1, ack => convTranspose_CP_39_elements(389)); -- 
    req_2984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(389), ack => WPIPE_Block3_start_1187_inst_req_0); -- 
    -- CP-element group 390:  transition  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (6) 
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_Update/req
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_Sample/ack
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_update_start_
      -- 
    ack_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1187_inst_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    req_2989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => WPIPE_Block3_start_1187_inst_req_1); -- 
    -- CP-element group 391:  transition  input  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (6) 
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_Sample/req
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_Sample/$entry
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_sample_start_
      -- CP-element group 391: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1187_Update/ack
      -- 
    ack_2990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1187_inst_ack_1, ack => convTranspose_CP_39_elements(391)); -- 
    req_2998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(391), ack => WPIPE_Block3_start_1190_inst_req_0); -- 
    -- CP-element group 392:  transition  input  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	393 
    -- CP-element group 392:  members (6) 
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_Update/req
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_Update/$entry
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_Sample/ack
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_update_start_
      -- CP-element group 392: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_sample_completed_
      -- 
    ack_2999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1190_inst_ack_0, ack => convTranspose_CP_39_elements(392)); -- 
    req_3003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(392), ack => WPIPE_Block3_start_1190_inst_req_1); -- 
    -- CP-element group 393:  transition  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	392 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (6) 
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_Sample/req
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_Update/ack
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1190_update_completed_
      -- 
    ack_3004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1190_inst_ack_1, ack => convTranspose_CP_39_elements(393)); -- 
    req_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(393), ack => WPIPE_Block3_start_1193_inst_req_0); -- 
    -- CP-element group 394:  transition  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (6) 
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_Update/req
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_Sample/ack
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_update_start_
      -- CP-element group 394: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_sample_completed_
      -- 
    ack_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1193_inst_ack_0, ack => convTranspose_CP_39_elements(394)); -- 
    req_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(394), ack => WPIPE_Block3_start_1193_inst_req_1); -- 
    -- CP-element group 395:  transition  input  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (6) 
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_Sample/req
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_Sample/$entry
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_sample_start_
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_Update/ack
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1193_update_completed_
      -- 
    ack_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1193_inst_ack_1, ack => convTranspose_CP_39_elements(395)); -- 
    req_3026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(395), ack => WPIPE_Block3_start_1196_inst_req_0); -- 
    -- CP-element group 396:  transition  input  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (6) 
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_Update/req
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_Update/$entry
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_Sample/ack
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_update_start_
      -- CP-element group 396: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_sample_completed_
      -- 
    ack_3027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1196_inst_ack_0, ack => convTranspose_CP_39_elements(396)); -- 
    req_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(396), ack => WPIPE_Block3_start_1196_inst_req_1); -- 
    -- CP-element group 397:  transition  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (6) 
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_Sample/req
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_Update/ack
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1196_update_completed_
      -- 
    ack_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1196_inst_ack_1, ack => convTranspose_CP_39_elements(397)); -- 
    req_3040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => WPIPE_Block3_start_1199_inst_req_0); -- 
    -- CP-element group 398:  transition  input  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (6) 
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_Sample/$exit
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_update_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_Sample/ack
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_Update/req
      -- 
    ack_3041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1199_inst_ack_0, ack => convTranspose_CP_39_elements(398)); -- 
    req_3045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => WPIPE_Block3_start_1199_inst_req_1); -- 
    -- CP-element group 399:  transition  input  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (6) 
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_Update/$exit
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1199_Update/ack
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_sample_start_
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_Sample/$entry
      -- 
    ack_3046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1199_inst_ack_1, ack => convTranspose_CP_39_elements(399)); -- 
    req_3054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(399), ack => WPIPE_Block3_start_1202_inst_req_0); -- 
    -- CP-element group 400:  transition  input  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (6) 
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_update_start_
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_sample_completed_
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_Update/req
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_Sample/ack
      -- CP-element group 400: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_Sample/$exit
      -- 
    ack_3055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1202_inst_ack_0, ack => convTranspose_CP_39_elements(400)); -- 
    req_3059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(400), ack => WPIPE_Block3_start_1202_inst_req_1); -- 
    -- CP-element group 401:  transition  input  output  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (6) 
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_update_completed_
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_Sample/req
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_Update/ack
      -- CP-element group 401: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1202_Update/$exit
      -- 
    ack_3060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1202_inst_ack_1, ack => convTranspose_CP_39_elements(401)); -- 
    req_3068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(401), ack => WPIPE_Block3_start_1205_inst_req_0); -- 
    -- CP-element group 402:  transition  input  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (6) 
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_Update/req
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_Sample/ack
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_Sample/$exit
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_update_start_
      -- CP-element group 402: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_sample_completed_
      -- 
    ack_3069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1205_inst_ack_0, ack => convTranspose_CP_39_elements(402)); -- 
    req_3073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => WPIPE_Block3_start_1205_inst_req_1); -- 
    -- CP-element group 403:  transition  input  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (6) 
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_Sample/req
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_Sample/$entry
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_sample_start_
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_Update/ack
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_Update/$exit
      -- CP-element group 403: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1205_update_completed_
      -- 
    ack_3074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1205_inst_ack_1, ack => convTranspose_CP_39_elements(403)); -- 
    req_3082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(403), ack => WPIPE_Block3_start_1208_inst_req_0); -- 
    -- CP-element group 404:  transition  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (6) 
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_Update/req
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_Sample/ack
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_Sample/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_sample_completed_
      -- 
    ack_3083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1208_inst_ack_0, ack => convTranspose_CP_39_elements(404)); -- 
    req_3087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => WPIPE_Block3_start_1208_inst_req_1); -- 
    -- CP-element group 405:  transition  input  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (6) 
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_Sample/req
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_sample_start_
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_Update/ack
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1208_update_completed_
      -- 
    ack_3088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1208_inst_ack_1, ack => convTranspose_CP_39_elements(405)); -- 
    req_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(405), ack => WPIPE_Block3_start_1211_inst_req_0); -- 
    -- CP-element group 406:  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (6) 
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_Update/req
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_Sample/ack
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_Sample/$exit
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_update_start_
      -- CP-element group 406: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_sample_completed_
      -- 
    ack_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1211_inst_ack_0, ack => convTranspose_CP_39_elements(406)); -- 
    req_3101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(406), ack => WPIPE_Block3_start_1211_inst_req_1); -- 
    -- CP-element group 407:  transition  input  output  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (6) 
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_Sample/req
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_Sample/$entry
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_sample_start_
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_Update/ack
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_Update/$exit
      -- CP-element group 407: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1211_update_completed_
      -- 
    ack_3102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1211_inst_ack_1, ack => convTranspose_CP_39_elements(407)); -- 
    req_3110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(407), ack => WPIPE_Block3_start_1214_inst_req_0); -- 
    -- CP-element group 408:  transition  input  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (6) 
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_Sample/ack
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_Update/$entry
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_Update/req
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_Sample/$exit
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_update_start_
      -- CP-element group 408: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_sample_completed_
      -- 
    ack_3111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1214_inst_ack_0, ack => convTranspose_CP_39_elements(408)); -- 
    req_3115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(408), ack => WPIPE_Block3_start_1214_inst_req_1); -- 
    -- CP-element group 409:  transition  input  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (6) 
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_Sample/$entry
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_sample_start_
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_Update/ack
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_Update/$exit
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_Sample/req
      -- CP-element group 409: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1214_update_completed_
      -- 
    ack_3116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1214_inst_ack_1, ack => convTranspose_CP_39_elements(409)); -- 
    req_3124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(409), ack => WPIPE_Block3_start_1217_inst_req_0); -- 
    -- CP-element group 410:  transition  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (6) 
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_Sample/ack
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_Update/req
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_update_start_
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_Sample/$exit
      -- CP-element group 410: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_Update/$entry
      -- 
    ack_3125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1217_inst_ack_0, ack => convTranspose_CP_39_elements(410)); -- 
    req_3129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(410), ack => WPIPE_Block3_start_1217_inst_req_1); -- 
    -- CP-element group 411:  transition  input  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (6) 
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_Update/ack
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_Update/$exit
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1217_update_completed_
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_Sample/req
      -- CP-element group 411: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_Sample/$entry
      -- 
    ack_3130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1217_inst_ack_1, ack => convTranspose_CP_39_elements(411)); -- 
    req_3138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(411), ack => WPIPE_Block3_start_1220_inst_req_0); -- 
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_Update/req
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_Sample/ack
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_update_start_
      -- 
    ack_3139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1220_inst_ack_0, ack => convTranspose_CP_39_elements(412)); -- 
    req_3143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(412), ack => WPIPE_Block3_start_1220_inst_req_1); -- 
    -- CP-element group 413:  transition  input  output  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (6) 
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_Sample/req
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_Sample/$entry
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_sample_start_
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_Update/ack
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1220_update_completed_
      -- 
    ack_3144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1220_inst_ack_1, ack => convTranspose_CP_39_elements(413)); -- 
    req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(413), ack => WPIPE_Block3_start_1223_inst_req_0); -- 
    -- CP-element group 414:  transition  input  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (6) 
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_Update/req
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_Sample/ack
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_Sample/$exit
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_update_start_
      -- CP-element group 414: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_sample_completed_
      -- 
    ack_3153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 414_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1223_inst_ack_0, ack => convTranspose_CP_39_elements(414)); -- 
    req_3157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(414), ack => WPIPE_Block3_start_1223_inst_req_1); -- 
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_Sample/req
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_Sample/$entry
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_sample_start_
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_Update/ack
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_Update/$exit
      -- CP-element group 415: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1223_update_completed_
      -- 
    ack_3158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1223_inst_ack_1, ack => convTranspose_CP_39_elements(415)); -- 
    req_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(415), ack => WPIPE_Block3_start_1226_inst_req_0); -- 
    -- CP-element group 416:  transition  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416:  members (6) 
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_Update/req
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_Update/$entry
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_Sample/ack
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_update_start_
      -- CP-element group 416: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_sample_completed_
      -- 
    ack_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1226_inst_ack_0, ack => convTranspose_CP_39_elements(416)); -- 
    req_3171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(416), ack => WPIPE_Block3_start_1226_inst_req_1); -- 
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	420 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_Update/ack
      -- CP-element group 417: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1226_update_completed_
      -- 
    ack_3172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1226_inst_ack_1, ack => convTranspose_CP_39_elements(417)); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	528 
    -- CP-element group 418: successors 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_Sample/ra
      -- CP-element group 418: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_Sample/$exit
      -- CP-element group 418: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_sample_completed_
      -- 
    ra_3181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => convTranspose_CP_39_elements(418)); -- 
    -- CP-element group 419:  fork  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	528 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	420 
    -- CP-element group 419: 	423 
    -- CP-element group 419: 	426 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_Update/ca
      -- CP-element group 419: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_Update/$exit
      -- CP-element group 419: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_update_completed_
      -- 
    ca_3186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => convTranspose_CP_39_elements(419)); -- 
    -- CP-element group 420:  join  transition  output  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	417 
    -- CP-element group 420: 	419 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	421 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_Sample/req
      -- CP-element group 420: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_Sample/$entry
      -- CP-element group 420: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_sample_start_
      -- 
    req_3194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(420), ack => WPIPE_Block3_start_1240_inst_req_0); -- 
    convTranspose_cp_element_group_420: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_420"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(417) & convTranspose_CP_39_elements(419);
      gj_convTranspose_cp_element_group_420 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(420), clk => clk, reset => reset); --
    end block;
    -- CP-element group 421:  transition  input  output  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	420 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (6) 
      -- CP-element group 421: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_Update/req
      -- CP-element group 421: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_Update/$entry
      -- CP-element group 421: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_Sample/ack
      -- CP-element group 421: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_Sample/$exit
      -- CP-element group 421: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_update_start_
      -- CP-element group 421: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_sample_completed_
      -- 
    ack_3195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1240_inst_ack_0, ack => convTranspose_CP_39_elements(421)); -- 
    req_3199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(421), ack => WPIPE_Block3_start_1240_inst_req_1); -- 
    -- CP-element group 422:  transition  input  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_Update/ack
      -- CP-element group 422: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_Update/$exit
      -- CP-element group 422: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1240_update_completed_
      -- 
    ack_3200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1240_inst_ack_1, ack => convTranspose_CP_39_elements(422)); -- 
    -- CP-element group 423:  join  transition  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	419 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	424 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_Sample/req
      -- CP-element group 423: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_Sample/$entry
      -- CP-element group 423: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_sample_start_
      -- 
    req_3208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(423), ack => WPIPE_Block3_start_1243_inst_req_0); -- 
    convTranspose_cp_element_group_423: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_423"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(419) & convTranspose_CP_39_elements(422);
      gj_convTranspose_cp_element_group_423 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 424:  transition  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	423 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (6) 
      -- CP-element group 424: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_sample_completed_
      -- CP-element group 424: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_Sample/$exit
      -- CP-element group 424: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_Sample/ack
      -- CP-element group 424: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_Update/req
      -- CP-element group 424: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_update_start_
      -- 
    ack_3209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1243_inst_ack_0, ack => convTranspose_CP_39_elements(424)); -- 
    req_3213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(424), ack => WPIPE_Block3_start_1243_inst_req_1); -- 
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	426 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_Update/$exit
      -- CP-element group 425: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_Update/ack
      -- CP-element group 425: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1243_update_completed_
      -- 
    ack_3214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1243_inst_ack_1, ack => convTranspose_CP_39_elements(425)); -- 
    -- CP-element group 426:  join  transition  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	419 
    -- CP-element group 426: 	425 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_Sample/req
      -- 
    req_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(426), ack => WPIPE_Block3_start_1246_inst_req_0); -- 
    convTranspose_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(419) & convTranspose_CP_39_elements(425);
      gj_convTranspose_cp_element_group_426 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  transition  input  output  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (6) 
      -- CP-element group 427: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_sample_completed_
      -- CP-element group 427: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_update_start_
      -- CP-element group 427: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_Sample/$exit
      -- CP-element group 427: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_Sample/ack
      -- CP-element group 427: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_Update/req
      -- 
    ack_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1246_inst_ack_0, ack => convTranspose_CP_39_elements(427)); -- 
    req_3227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(427), ack => WPIPE_Block3_start_1246_inst_req_1); -- 
    -- CP-element group 428:  transition  input  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (6) 
      -- CP-element group 428: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_update_completed_
      -- CP-element group 428: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_Sample/req
      -- CP-element group 428: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_Sample/$entry
      -- CP-element group 428: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_sample_start_
      -- CP-element group 428: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_Update/ack
      -- CP-element group 428: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1246_Update/$exit
      -- 
    ack_3228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1246_inst_ack_1, ack => convTranspose_CP_39_elements(428)); -- 
    req_3236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(428), ack => WPIPE_Block3_start_1249_inst_req_0); -- 
    -- CP-element group 429:  transition  input  output  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (6) 
      -- CP-element group 429: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_Update/req
      -- CP-element group 429: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_Update/$entry
      -- CP-element group 429: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_Sample/ack
      -- CP-element group 429: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_Sample/$exit
      -- CP-element group 429: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_update_start_
      -- CP-element group 429: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_sample_completed_
      -- 
    ack_3237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1249_inst_ack_0, ack => convTranspose_CP_39_elements(429)); -- 
    req_3241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(429), ack => WPIPE_Block3_start_1249_inst_req_1); -- 
    -- CP-element group 430:  transition  input  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	431 
    -- CP-element group 430:  members (6) 
      -- CP-element group 430: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_Sample/req
      -- CP-element group 430: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_Update/ack
      -- CP-element group 430: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_Update/$exit
      -- CP-element group 430: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1249_update_completed_
      -- 
    ack_3242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1249_inst_ack_1, ack => convTranspose_CP_39_elements(430)); -- 
    req_3250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(430), ack => WPIPE_Block3_start_1252_inst_req_0); -- 
    -- CP-element group 431:  transition  input  output  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	430 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	432 
    -- CP-element group 431:  members (6) 
      -- CP-element group 431: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_Update/req
      -- CP-element group 431: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_Update/$entry
      -- CP-element group 431: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_Sample/ack
      -- CP-element group 431: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_update_start_
      -- CP-element group 431: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_sample_completed_
      -- 
    ack_3251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1252_inst_ack_0, ack => convTranspose_CP_39_elements(431)); -- 
    req_3255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(431), ack => WPIPE_Block3_start_1252_inst_req_1); -- 
    -- CP-element group 432:  transition  input  output  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	431 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	433 
    -- CP-element group 432:  members (6) 
      -- CP-element group 432: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_Sample/$entry
      -- CP-element group 432: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_sample_start_
      -- CP-element group 432: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_Update/ack
      -- CP-element group 432: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_Sample/req
      -- CP-element group 432: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1252_update_completed_
      -- 
    ack_3256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1252_inst_ack_1, ack => convTranspose_CP_39_elements(432)); -- 
    req_3264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(432), ack => WPIPE_Block3_start_1255_inst_req_0); -- 
    -- CP-element group 433:  transition  input  output  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	432 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	434 
    -- CP-element group 433:  members (6) 
      -- CP-element group 433: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_Update/$entry
      -- CP-element group 433: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_Sample/ack
      -- CP-element group 433: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_update_start_
      -- CP-element group 433: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_Update/req
      -- CP-element group 433: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_sample_completed_
      -- CP-element group 433: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_Sample/$exit
      -- 
    ack_3265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1255_inst_ack_0, ack => convTranspose_CP_39_elements(433)); -- 
    req_3269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(433), ack => WPIPE_Block3_start_1255_inst_req_1); -- 
    -- CP-element group 434:  transition  input  output  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	433 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	435 
    -- CP-element group 434:  members (6) 
      -- CP-element group 434: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_Update/$exit
      -- CP-element group 434: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_Update/ack
      -- CP-element group 434: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1255_update_completed_
      -- CP-element group 434: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_sample_start_
      -- CP-element group 434: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_Sample/req
      -- CP-element group 434: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_Sample/$entry
      -- 
    ack_3270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1255_inst_ack_1, ack => convTranspose_CP_39_elements(434)); -- 
    req_3278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(434), ack => WPIPE_Block3_start_1258_inst_req_0); -- 
    -- CP-element group 435:  transition  input  output  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	434 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	436 
    -- CP-element group 435:  members (6) 
      -- CP-element group 435: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_Update/req
      -- CP-element group 435: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_Update/$entry
      -- CP-element group 435: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_Sample/ack
      -- CP-element group 435: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_update_start_
      -- CP-element group 435: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_sample_completed_
      -- 
    ack_3279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1258_inst_ack_0, ack => convTranspose_CP_39_elements(435)); -- 
    req_3283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(435), ack => WPIPE_Block3_start_1258_inst_req_1); -- 
    -- CP-element group 436:  transition  input  output  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	435 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	437 
    -- CP-element group 436:  members (6) 
      -- CP-element group 436: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_Sample/req
      -- CP-element group 436: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_Sample/$entry
      -- CP-element group 436: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_sample_start_
      -- CP-element group 436: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_Update/ack
      -- CP-element group 436: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_Update/$exit
      -- CP-element group 436: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1258_update_completed_
      -- 
    ack_3284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1258_inst_ack_1, ack => convTranspose_CP_39_elements(436)); -- 
    req_3292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(436), ack => WPIPE_Block3_start_1261_inst_req_0); -- 
    -- CP-element group 437:  transition  input  output  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	436 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	438 
    -- CP-element group 437:  members (6) 
      -- CP-element group 437: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_Update/req
      -- CP-element group 437: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_Update/$entry
      -- CP-element group 437: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_Sample/ack
      -- CP-element group 437: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_Sample/$exit
      -- CP-element group 437: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_update_start_
      -- CP-element group 437: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_sample_completed_
      -- 
    ack_3293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1261_inst_ack_0, ack => convTranspose_CP_39_elements(437)); -- 
    req_3297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(437), ack => WPIPE_Block3_start_1261_inst_req_1); -- 
    -- CP-element group 438:  transition  input  output  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	437 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	439 
    -- CP-element group 438:  members (6) 
      -- CP-element group 438: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_sample_start_
      -- CP-element group 438: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_Update/ack
      -- CP-element group 438: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_Sample/$entry
      -- CP-element group 438: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_Update/$exit
      -- CP-element group 438: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1261_update_completed_
      -- CP-element group 438: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_Sample/req
      -- 
    ack_3298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1261_inst_ack_1, ack => convTranspose_CP_39_elements(438)); -- 
    req_3306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(438), ack => WPIPE_Block3_start_1264_inst_req_0); -- 
    -- CP-element group 439:  transition  input  output  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	438 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	440 
    -- CP-element group 439:  members (6) 
      -- CP-element group 439: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_sample_completed_
      -- CP-element group 439: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_update_start_
      -- CP-element group 439: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_Update/$entry
      -- CP-element group 439: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_Update/req
      -- CP-element group 439: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_Sample/ack
      -- CP-element group 439: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_Sample/$exit
      -- 
    ack_3307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1264_inst_ack_0, ack => convTranspose_CP_39_elements(439)); -- 
    req_3311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(439), ack => WPIPE_Block3_start_1264_inst_req_1); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	439 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	449 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_Update/ack
      -- CP-element group 440: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_Update/$exit
      -- CP-element group 440: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1264_update_completed_
      -- 
    ack_3312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1264_inst_ack_1, ack => convTranspose_CP_39_elements(440)); -- 
    -- CP-element group 441:  transition  input  output  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	528 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441:  members (6) 
      -- CP-element group 441: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_Sample/$exit
      -- CP-element group 441: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_Update/$entry
      -- CP-element group 441: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_sample_completed_
      -- CP-element group 441: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_update_start_
      -- CP-element group 441: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_Sample/ra
      -- CP-element group 441: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_Update/cr
      -- 
    ra_3321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1268_inst_ack_0, ack => convTranspose_CP_39_elements(441)); -- 
    cr_3325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(441), ack => RPIPE_Block0_done_1268_inst_req_1); -- 
    -- CP-element group 442:  transition  input  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	441 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	449 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_Update/$exit
      -- CP-element group 442: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_update_completed_
      -- CP-element group 442: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_Update/ca
      -- 
    ca_3326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1268_inst_ack_1, ack => convTranspose_CP_39_elements(442)); -- 
    -- CP-element group 443:  transition  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	528 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (6) 
      -- CP-element group 443: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_Sample/ra
      -- CP-element group 443: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_update_start_
      -- CP-element group 443: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_sample_completed_
      -- 
    ra_3335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1271_inst_ack_0, ack => convTranspose_CP_39_elements(443)); -- 
    cr_3339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(443), ack => RPIPE_Block1_done_1271_inst_req_1); -- 
    -- CP-element group 444:  transition  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	449 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_Update/ca
      -- CP-element group 444: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_update_completed_
      -- 
    ca_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1271_inst_ack_1, ack => convTranspose_CP_39_elements(444)); -- 
    -- CP-element group 445:  transition  input  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	528 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (6) 
      -- CP-element group 445: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_Update/cr
      -- CP-element group 445: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_Update/$entry
      -- CP-element group 445: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_Sample/ra
      -- CP-element group 445: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_Sample/$exit
      -- CP-element group 445: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_update_start_
      -- CP-element group 445: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_sample_completed_
      -- 
    ra_3349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1274_inst_ack_0, ack => convTranspose_CP_39_elements(445)); -- 
    cr_3353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(445), ack => RPIPE_Block2_done_1274_inst_req_1); -- 
    -- CP-element group 446:  transition  input  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	449 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_Update/ca
      -- CP-element group 446: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_Update/$exit
      -- CP-element group 446: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_update_completed_
      -- 
    ca_3354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1274_inst_ack_1, ack => convTranspose_CP_39_elements(446)); -- 
    -- CP-element group 447:  transition  input  output  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	528 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (6) 
      -- CP-element group 447: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_sample_completed_
      -- CP-element group 447: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_update_start_
      -- CP-element group 447: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_Sample/$exit
      -- CP-element group 447: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_Sample/ra
      -- CP-element group 447: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_Update/$entry
      -- CP-element group 447: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_Update/cr
      -- 
    ra_3363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1277_inst_ack_0, ack => convTranspose_CP_39_elements(447)); -- 
    cr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(447), ack => RPIPE_Block3_done_1277_inst_req_1); -- 
    -- CP-element group 448:  transition  input  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_update_completed_
      -- CP-element group 448: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_Update/ca
      -- CP-element group 448: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_Update/$exit
      -- 
    ca_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1277_inst_ack_1, ack => convTranspose_CP_39_elements(448)); -- 
    -- CP-element group 449:  join  fork  transition  place  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	198 
    -- CP-element group 449: 	254 
    -- CP-element group 449: 	318 
    -- CP-element group 449: 	379 
    -- CP-element group 449: 	440 
    -- CP-element group 449: 	442 
    -- CP-element group 449: 	444 
    -- CP-element group 449: 	446 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449: 	451 
    -- CP-element group 449: 	453 
    -- CP-element group 449:  members (13) 
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278__exit__
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294__entry__
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/$exit
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_sample_start_
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_update_start_
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_Sample/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_Sample/crr
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_Update/ccr
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_update_start_
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_Update/cr
      -- 
    crr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(449), ack => call_stmt_1281_call_req_0); -- 
    ccr_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(449), ack => call_stmt_1281_call_req_1); -- 
    cr_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(449), ack => type_cast_1285_inst_req_1); -- 
    convTranspose_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(198) & convTranspose_CP_39_elements(254) & convTranspose_CP_39_elements(318) & convTranspose_CP_39_elements(379) & convTranspose_CP_39_elements(440) & convTranspose_CP_39_elements(442) & convTranspose_CP_39_elements(444) & convTranspose_CP_39_elements(446) & convTranspose_CP_39_elements(448);
      gj_convTranspose_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  transition  input  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_sample_completed_
      -- CP-element group 450: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_Sample/$exit
      -- CP-element group 450: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_Sample/cra
      -- 
    cra_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1281_call_ack_0, ack => convTranspose_CP_39_elements(450)); -- 
    -- CP-element group 451:  transition  input  output  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	449 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (6) 
      -- CP-element group 451: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_update_completed_
      -- CP-element group 451: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_Update/$exit
      -- CP-element group 451: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/call_stmt_1281_Update/cca
      -- CP-element group 451: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_sample_start_
      -- CP-element group 451: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_Sample/rr
      -- 
    cca_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1281_call_ack_1, ack => convTranspose_CP_39_elements(451)); -- 
    rr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(451), ack => type_cast_1285_inst_req_0); -- 
    -- CP-element group 452:  transition  input  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_sample_completed_
      -- CP-element group 452: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_Sample/ra
      -- 
    ra_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1285_inst_ack_0, ack => convTranspose_CP_39_elements(452)); -- 
    -- CP-element group 453:  transition  input  output  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	449 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (6) 
      -- CP-element group 453: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_update_completed_
      -- CP-element group 453: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/type_cast_1285_Update/ca
      -- CP-element group 453: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_sample_start_
      -- CP-element group 453: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_Sample/$entry
      -- CP-element group 453: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_Sample/req
      -- 
    ca_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1285_inst_ack_1, ack => convTranspose_CP_39_elements(453)); -- 
    req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(453), ack => WPIPE_elapsed_time_pipe_1292_inst_req_0); -- 
    -- CP-element group 454:  transition  input  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (6) 
      -- CP-element group 454: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_sample_completed_
      -- CP-element group 454: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_update_start_
      -- CP-element group 454: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_Sample/$exit
      -- CP-element group 454: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_Sample/ack
      -- CP-element group 454: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_Update/$entry
      -- CP-element group 454: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_Update/req
      -- 
    ack_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 454_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1292_inst_ack_0, ack => convTranspose_CP_39_elements(454)); -- 
    req_3412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(454), ack => WPIPE_elapsed_time_pipe_1292_inst_req_1); -- 
    -- CP-element group 455:  branch  transition  place  input  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455: 	457 
    -- CP-element group 455:  members (13) 
      -- CP-element group 455: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294__exit__
      -- CP-element group 455: 	 branch_block_stmt_32/if_stmt_1296__entry__
      -- CP-element group 455: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/$exit
      -- CP-element group 455: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_update_completed_
      -- CP-element group 455: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_Update/$exit
      -- CP-element group 455: 	 branch_block_stmt_32/call_stmt_1281_to_assign_stmt_1294/WPIPE_elapsed_time_pipe_1292_Update/ack
      -- CP-element group 455: 	 branch_block_stmt_32/if_stmt_1296_dead_link/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/if_stmt_1296_eval_test/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/if_stmt_1296_eval_test/$exit
      -- CP-element group 455: 	 branch_block_stmt_32/if_stmt_1296_eval_test/branch_req
      -- CP-element group 455: 	 branch_block_stmt_32/R_cmp264755_1297_place
      -- CP-element group 455: 	 branch_block_stmt_32/if_stmt_1296_if_link/$entry
      -- CP-element group 455: 	 branch_block_stmt_32/if_stmt_1296_else_link/$entry
      -- 
    ack_3413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1292_inst_ack_1, ack => convTranspose_CP_39_elements(455)); -- 
    branch_req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(455), ack => if_stmt_1296_branch_req_0); -- 
    -- CP-element group 456:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	458 
    -- CP-element group 456: 	459 
    -- CP-element group 456:  members (18) 
      -- CP-element group 456: 	 branch_block_stmt_32/merge_stmt_1302__exit__
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337__entry__
      -- CP-element group 456: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 456: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 456: 	 branch_block_stmt_32/merge_stmt_1302_PhiAck/$entry
      -- CP-element group 456: 	 branch_block_stmt_32/merge_stmt_1302_PhiAck/$exit
      -- CP-element group 456: 	 branch_block_stmt_32/merge_stmt_1302_PhiAck/dummy
      -- CP-element group 456: 	 branch_block_stmt_32/if_stmt_1296_if_link/$exit
      -- CP-element group 456: 	 branch_block_stmt_32/if_stmt_1296_if_link/if_choice_transition
      -- CP-element group 456: 	 branch_block_stmt_32/forx_xend273_bbx_xnph
      -- CP-element group 456: 	 branch_block_stmt_32/merge_stmt_1302_PhiReqMerge
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/$entry
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_sample_start_
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_update_start_
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_Sample/$entry
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_Sample/rr
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_Update/$entry
      -- CP-element group 456: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_Update/cr
      -- 
    if_choice_transition_3426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1296_branch_ack_1, ack => convTranspose_CP_39_elements(456)); -- 
    rr_3443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(456), ack => type_cast_1323_inst_req_0); -- 
    cr_3448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(456), ack => type_cast_1323_inst_req_1); -- 
    -- CP-element group 457:  transition  place  input  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	455 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	535 
    -- CP-element group 457:  members (5) 
      -- CP-element group 457: 	 branch_block_stmt_32/forx_xend273_forx_xend702_PhiReq/$entry
      -- CP-element group 457: 	 branch_block_stmt_32/forx_xend273_forx_xend702_PhiReq/$exit
      -- CP-element group 457: 	 branch_block_stmt_32/if_stmt_1296_else_link/$exit
      -- CP-element group 457: 	 branch_block_stmt_32/if_stmt_1296_else_link/else_choice_transition
      -- CP-element group 457: 	 branch_block_stmt_32/forx_xend273_forx_xend702
      -- 
    else_choice_transition_3430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1296_branch_ack_0, ack => convTranspose_CP_39_elements(457)); -- 
    -- CP-element group 458:  transition  input  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	456 
    -- CP-element group 458: successors 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_sample_completed_
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_Sample/$exit
      -- CP-element group 458: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_Sample/ra
      -- 
    ra_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1323_inst_ack_0, ack => convTranspose_CP_39_elements(458)); -- 
    -- CP-element group 459:  transition  place  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	456 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	529 
    -- CP-element group 459:  members (9) 
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337__exit__
      -- CP-element group 459: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630
      -- CP-element group 459: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630_PhiReq/$entry
      -- CP-element group 459: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630_PhiReq/phi_stmt_1340/$entry
      -- CP-element group 459: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/$entry
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_update_completed_
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_Update/$exit
      -- CP-element group 459: 	 branch_block_stmt_32/assign_stmt_1308_to_assign_stmt_1337/type_cast_1323_Update/ca
      -- 
    ca_3449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1323_inst_ack_1, ack => convTranspose_CP_39_elements(459)); -- 
    -- CP-element group 460:  transition  input  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	534 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	505 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_sample_complete
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_Sample/$exit
      -- CP-element group 460: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_Sample/ack
      -- 
    ack_3478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1352_index_offset_ack_0, ack => convTranspose_CP_39_elements(460)); -- 
    -- CP-element group 461:  transition  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	534 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (11) 
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_sample_start_
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_root_address_calculated
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_offset_calculated
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_Update/$exit
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_Update/ack
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_base_plus_offset/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_base_plus_offset/$exit
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_base_plus_offset/sum_rename_req
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_base_plus_offset/sum_rename_ack
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_request/$entry
      -- CP-element group 461: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_request/req
      -- 
    ack_3483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1352_index_offset_ack_1, ack => convTranspose_CP_39_elements(461)); -- 
    req_3492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(461), ack => addr_of_1353_final_reg_req_0); -- 
    -- CP-element group 462:  transition  input  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_sample_completed_
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_request/$exit
      -- CP-element group 462: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_request/ack
      -- 
    ack_3493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1353_final_reg_ack_0, ack => convTranspose_CP_39_elements(462)); -- 
    -- CP-element group 463:  join  fork  transition  input  output  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	534 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (24) 
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_update_completed_
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_complete/$exit
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_complete/ack
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_address_calculated
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_word_address_calculated
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_root_address_calculated
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_address_resized
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_addr_resize/$entry
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_addr_resize/$exit
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_addr_resize/base_resize_req
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_addr_resize/base_resize_ack
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_plus_offset/$entry
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_plus_offset/$exit
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_plus_offset/sum_rename_req
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_base_plus_offset/sum_rename_ack
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_word_addrgen/$entry
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_word_addrgen/$exit
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_word_addrgen/root_register_req
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_word_addrgen/root_register_ack
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Sample/$entry
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Sample/word_access_start/$entry
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Sample/word_access_start/word_0/$entry
      -- CP-element group 463: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Sample/word_access_start/word_0/rr
      -- 
    ack_3498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1353_final_reg_ack_1, ack => convTranspose_CP_39_elements(463)); -- 
    rr_3531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(463), ack => ptr_deref_1357_load_0_req_0); -- 
    -- CP-element group 464:  transition  input  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464:  members (5) 
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Sample/word_access_start/$exit
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Sample/word_access_start/word_0/$exit
      -- CP-element group 464: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Sample/word_access_start/word_0/ra
      -- 
    ra_3532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_load_0_ack_0, ack => convTranspose_CP_39_elements(464)); -- 
    -- CP-element group 465:  fork  transition  input  output  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	534 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	470 
    -- CP-element group 465: 	472 
    -- CP-element group 465: 	474 
    -- CP-element group 465: 	476 
    -- CP-element group 465: 	478 
    -- CP-element group 465: 	480 
    -- CP-element group 465: 	466 
    -- CP-element group 465: 	468 
    -- CP-element group 465:  members (33) 
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/word_access_complete/$exit
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/word_access_complete/word_0/$exit
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/word_access_complete/word_0/ca
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/ptr_deref_1357_Merge/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/ptr_deref_1357_Merge/$exit
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/ptr_deref_1357_Merge/merge_req
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/ptr_deref_1357_Merge/merge_ack
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_Sample/rr
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_Sample/rr
      -- 
    ca_3543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_load_0_ack_1, ack => convTranspose_CP_39_elements(465)); -- 
    rr_3584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(465), ack => type_cast_1381_inst_req_0); -- 
    rr_3598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(465), ack => type_cast_1391_inst_req_0); -- 
    rr_3612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(465), ack => type_cast_1401_inst_req_0); -- 
    rr_3626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(465), ack => type_cast_1411_inst_req_0); -- 
    rr_3640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(465), ack => type_cast_1421_inst_req_0); -- 
    rr_3654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(465), ack => type_cast_1431_inst_req_0); -- 
    rr_3556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(465), ack => type_cast_1361_inst_req_0); -- 
    rr_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(465), ack => type_cast_1371_inst_req_0); -- 
    -- CP-element group 466:  transition  input  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_sample_completed_
      -- CP-element group 466: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_Sample/$exit
      -- CP-element group 466: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_Sample/ra
      -- 
    ra_3557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 466_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_0, ack => convTranspose_CP_39_elements(466)); -- 
    -- CP-element group 467:  transition  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	534 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	502 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_update_completed_
      -- CP-element group 467: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_Update/$exit
      -- CP-element group 467: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_Update/ca
      -- 
    ca_3562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_1, ack => convTranspose_CP_39_elements(467)); -- 
    -- CP-element group 468:  transition  input  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	465 
    -- CP-element group 468: successors 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_sample_completed_
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_Sample/$exit
      -- CP-element group 468: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_Sample/ra
      -- 
    ra_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_0, ack => convTranspose_CP_39_elements(468)); -- 
    -- CP-element group 469:  transition  input  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	534 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	499 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_update_completed_
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_Update/$exit
      -- CP-element group 469: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_Update/ca
      -- 
    ca_3576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1371_inst_ack_1, ack => convTranspose_CP_39_elements(469)); -- 
    -- CP-element group 470:  transition  input  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	465 
    -- CP-element group 470: successors 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_sample_completed_
      -- CP-element group 470: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_Sample/$exit
      -- CP-element group 470: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_Sample/ra
      -- 
    ra_3585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 470_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1381_inst_ack_0, ack => convTranspose_CP_39_elements(470)); -- 
    -- CP-element group 471:  transition  input  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	534 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	496 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_update_completed_
      -- CP-element group 471: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_Update/$exit
      -- CP-element group 471: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_Update/ca
      -- 
    ca_3590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1381_inst_ack_1, ack => convTranspose_CP_39_elements(471)); -- 
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	465 
    -- CP-element group 472: successors 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_sample_completed_
      -- CP-element group 472: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_Sample/$exit
      -- CP-element group 472: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_Sample/ra
      -- 
    ra_3599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_0, ack => convTranspose_CP_39_elements(472)); -- 
    -- CP-element group 473:  transition  input  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	534 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	493 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_update_completed_
      -- CP-element group 473: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_Update/$exit
      -- CP-element group 473: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_Update/ca
      -- 
    ca_3604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_1, ack => convTranspose_CP_39_elements(473)); -- 
    -- CP-element group 474:  transition  input  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	465 
    -- CP-element group 474: successors 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_sample_completed_
      -- CP-element group 474: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_Sample/$exit
      -- CP-element group 474: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_Sample/ra
      -- 
    ra_3613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 474_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1401_inst_ack_0, ack => convTranspose_CP_39_elements(474)); -- 
    -- CP-element group 475:  transition  input  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	534 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	490 
    -- CP-element group 475:  members (3) 
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_update_completed_
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_Update/$exit
      -- CP-element group 475: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_Update/ca
      -- 
    ca_3618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1401_inst_ack_1, ack => convTranspose_CP_39_elements(475)); -- 
    -- CP-element group 476:  transition  input  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	465 
    -- CP-element group 476: successors 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_sample_completed_
      -- CP-element group 476: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_Sample/$exit
      -- CP-element group 476: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_Sample/ra
      -- 
    ra_3627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_0, ack => convTranspose_CP_39_elements(476)); -- 
    -- CP-element group 477:  transition  input  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	534 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	487 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_update_completed_
      -- CP-element group 477: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_Update/$exit
      -- CP-element group 477: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_Update/ca
      -- 
    ca_3632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1411_inst_ack_1, ack => convTranspose_CP_39_elements(477)); -- 
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	465 
    -- CP-element group 478: successors 
    -- CP-element group 478:  members (3) 
      -- CP-element group 478: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_sample_completed_
      -- CP-element group 478: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_Sample/$exit
      -- CP-element group 478: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_Sample/ra
      -- 
    ra_3641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1421_inst_ack_0, ack => convTranspose_CP_39_elements(478)); -- 
    -- CP-element group 479:  transition  input  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	534 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	484 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_update_completed_
      -- CP-element group 479: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_Update/$exit
      -- CP-element group 479: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_Update/ca
      -- 
    ca_3646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1421_inst_ack_1, ack => convTranspose_CP_39_elements(479)); -- 
    -- CP-element group 480:  transition  input  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	465 
    -- CP-element group 480: successors 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_sample_completed_
      -- CP-element group 480: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_Sample/$exit
      -- CP-element group 480: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_Sample/ra
      -- 
    ra_3655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1431_inst_ack_0, ack => convTranspose_CP_39_elements(480)); -- 
    -- CP-element group 481:  transition  input  output  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	534 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	482 
    -- CP-element group 481:  members (6) 
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_update_completed_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_Update/$exit
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_Update/ca
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_sample_start_
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_Sample/req
      -- 
    ca_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1431_inst_ack_1, ack => convTranspose_CP_39_elements(481)); -- 
    req_3668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(481), ack => WPIPE_ConvTranspose_output_pipe_1433_inst_req_0); -- 
    -- CP-element group 482:  transition  input  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	481 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	483 
    -- CP-element group 482:  members (6) 
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_sample_completed_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_update_start_
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_Sample/$exit
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_Sample/ack
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_Update/req
      -- 
    ack_3669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 482_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1433_inst_ack_0, ack => convTranspose_CP_39_elements(482)); -- 
    req_3673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(482), ack => WPIPE_ConvTranspose_output_pipe_1433_inst_req_1); -- 
    -- CP-element group 483:  transition  input  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	482 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	484 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_update_completed_
      -- CP-element group 483: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_Update/$exit
      -- CP-element group 483: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1433_Update/ack
      -- 
    ack_3674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1433_inst_ack_1, ack => convTranspose_CP_39_elements(483)); -- 
    -- CP-element group 484:  join  transition  output  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	479 
    -- CP-element group 484: 	483 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	485 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_sample_start_
      -- CP-element group 484: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_Sample/$entry
      -- CP-element group 484: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_Sample/req
      -- 
    req_3682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(484), ack => WPIPE_ConvTranspose_output_pipe_1436_inst_req_0); -- 
    convTranspose_cp_element_group_484: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_484"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(479) & convTranspose_CP_39_elements(483);
      gj_convTranspose_cp_element_group_484 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(484), clk => clk, reset => reset); --
    end block;
    -- CP-element group 485:  transition  input  output  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	484 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	486 
    -- CP-element group 485:  members (6) 
      -- CP-element group 485: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_sample_completed_
      -- CP-element group 485: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_update_start_
      -- CP-element group 485: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_Sample/$exit
      -- CP-element group 485: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_Sample/ack
      -- CP-element group 485: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_Update/$entry
      -- CP-element group 485: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_Update/req
      -- 
    ack_3683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1436_inst_ack_0, ack => convTranspose_CP_39_elements(485)); -- 
    req_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(485), ack => WPIPE_ConvTranspose_output_pipe_1436_inst_req_1); -- 
    -- CP-element group 486:  transition  input  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	485 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_update_completed_
      -- CP-element group 486: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_Update/$exit
      -- CP-element group 486: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1436_Update/ack
      -- 
    ack_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 486_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1436_inst_ack_1, ack => convTranspose_CP_39_elements(486)); -- 
    -- CP-element group 487:  join  transition  output  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	477 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_sample_start_
      -- CP-element group 487: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_Sample/$entry
      -- CP-element group 487: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_Sample/req
      -- 
    req_3696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(487), ack => WPIPE_ConvTranspose_output_pipe_1439_inst_req_0); -- 
    convTranspose_cp_element_group_487: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_487"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(477) & convTranspose_CP_39_elements(486);
      gj_convTranspose_cp_element_group_487 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(487), clk => clk, reset => reset); --
    end block;
    -- CP-element group 488:  transition  input  output  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	489 
    -- CP-element group 488:  members (6) 
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_sample_completed_
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_update_start_
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_Sample/$exit
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_Sample/ack
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_Update/$entry
      -- CP-element group 488: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_Update/req
      -- 
    ack_3697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1439_inst_ack_0, ack => convTranspose_CP_39_elements(488)); -- 
    req_3701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(488), ack => WPIPE_ConvTranspose_output_pipe_1439_inst_req_1); -- 
    -- CP-element group 489:  transition  input  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	488 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	490 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_update_completed_
      -- CP-element group 489: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_Update/$exit
      -- CP-element group 489: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1439_Update/ack
      -- 
    ack_3702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1439_inst_ack_1, ack => convTranspose_CP_39_elements(489)); -- 
    -- CP-element group 490:  join  transition  output  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	475 
    -- CP-element group 490: 	489 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	491 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_sample_start_
      -- CP-element group 490: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_Sample/$entry
      -- CP-element group 490: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_Sample/req
      -- 
    req_3710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(490), ack => WPIPE_ConvTranspose_output_pipe_1442_inst_req_0); -- 
    convTranspose_cp_element_group_490: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_490"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(475) & convTranspose_CP_39_elements(489);
      gj_convTranspose_cp_element_group_490 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(490), clk => clk, reset => reset); --
    end block;
    -- CP-element group 491:  transition  input  output  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	490 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	492 
    -- CP-element group 491:  members (6) 
      -- CP-element group 491: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_sample_completed_
      -- CP-element group 491: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_update_start_
      -- CP-element group 491: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_Sample/ack
      -- CP-element group 491: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_Update/$entry
      -- CP-element group 491: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_Update/req
      -- 
    ack_3711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0, ack => convTranspose_CP_39_elements(491)); -- 
    req_3715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(491), ack => WPIPE_ConvTranspose_output_pipe_1442_inst_req_1); -- 
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	491 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492:  members (3) 
      -- CP-element group 492: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_update_completed_
      -- CP-element group 492: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1442_Update/ack
      -- 
    ack_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1, ack => convTranspose_CP_39_elements(492)); -- 
    -- CP-element group 493:  join  transition  output  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	473 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_sample_start_
      -- CP-element group 493: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_Sample/$entry
      -- CP-element group 493: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_Sample/req
      -- 
    req_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(493), ack => WPIPE_ConvTranspose_output_pipe_1445_inst_req_0); -- 
    convTranspose_cp_element_group_493: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_493"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(473) & convTranspose_CP_39_elements(492);
      gj_convTranspose_cp_element_group_493 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(493), clk => clk, reset => reset); --
    end block;
    -- CP-element group 494:  transition  input  output  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	493 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (6) 
      -- CP-element group 494: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_sample_completed_
      -- CP-element group 494: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_update_start_
      -- CP-element group 494: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_Sample/$exit
      -- CP-element group 494: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_Sample/ack
      -- CP-element group 494: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_Update/$entry
      -- CP-element group 494: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_Update/req
      -- 
    ack_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0, ack => convTranspose_CP_39_elements(494)); -- 
    req_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(494), ack => WPIPE_ConvTranspose_output_pipe_1445_inst_req_1); -- 
    -- CP-element group 495:  transition  input  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	496 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_update_completed_
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_Update/$exit
      -- CP-element group 495: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1445_Update/ack
      -- 
    ack_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1, ack => convTranspose_CP_39_elements(495)); -- 
    -- CP-element group 496:  join  transition  output  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	471 
    -- CP-element group 496: 	495 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	497 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_sample_start_
      -- CP-element group 496: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_Sample/$entry
      -- CP-element group 496: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_Sample/req
      -- 
    req_3738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(496), ack => WPIPE_ConvTranspose_output_pipe_1448_inst_req_0); -- 
    convTranspose_cp_element_group_496: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_496"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(471) & convTranspose_CP_39_elements(495);
      gj_convTranspose_cp_element_group_496 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(496), clk => clk, reset => reset); --
    end block;
    -- CP-element group 497:  transition  input  output  bypass 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	496 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	498 
    -- CP-element group 497:  members (6) 
      -- CP-element group 497: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_sample_completed_
      -- CP-element group 497: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_update_start_
      -- CP-element group 497: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_Sample/$exit
      -- CP-element group 497: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_Sample/ack
      -- CP-element group 497: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_Update/$entry
      -- CP-element group 497: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_Update/req
      -- 
    ack_3739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 497_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0, ack => convTranspose_CP_39_elements(497)); -- 
    req_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(497), ack => WPIPE_ConvTranspose_output_pipe_1448_inst_req_1); -- 
    -- CP-element group 498:  transition  input  bypass 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	497 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	499 
    -- CP-element group 498:  members (3) 
      -- CP-element group 498: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_update_completed_
      -- CP-element group 498: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_Update/$exit
      -- CP-element group 498: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1448_Update/ack
      -- 
    ack_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1, ack => convTranspose_CP_39_elements(498)); -- 
    -- CP-element group 499:  join  transition  output  bypass 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	498 
    -- CP-element group 499: 	469 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	500 
    -- CP-element group 499:  members (3) 
      -- CP-element group 499: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_sample_start_
      -- CP-element group 499: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_Sample/$entry
      -- CP-element group 499: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_Sample/req
      -- 
    req_3752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(499), ack => WPIPE_ConvTranspose_output_pipe_1451_inst_req_0); -- 
    convTranspose_cp_element_group_499: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_499"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(498) & convTranspose_CP_39_elements(469);
      gj_convTranspose_cp_element_group_499 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(499), clk => clk, reset => reset); --
    end block;
    -- CP-element group 500:  transition  input  output  bypass 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	499 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	501 
    -- CP-element group 500:  members (6) 
      -- CP-element group 500: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_sample_completed_
      -- CP-element group 500: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_update_start_
      -- CP-element group 500: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_Sample/$exit
      -- CP-element group 500: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_Sample/ack
      -- CP-element group 500: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_Update/$entry
      -- CP-element group 500: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_Update/req
      -- 
    ack_3753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0, ack => convTranspose_CP_39_elements(500)); -- 
    req_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(500), ack => WPIPE_ConvTranspose_output_pipe_1451_inst_req_1); -- 
    -- CP-element group 501:  transition  input  bypass 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	500 
    -- CP-element group 501: successors 
    -- CP-element group 501: 	502 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_update_completed_
      -- CP-element group 501: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_Update/$exit
      -- CP-element group 501: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1451_Update/ack
      -- 
    ack_3758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1, ack => convTranspose_CP_39_elements(501)); -- 
    -- CP-element group 502:  join  transition  output  bypass 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	501 
    -- CP-element group 502: 	467 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	503 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_sample_start_
      -- CP-element group 502: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_Sample/$entry
      -- CP-element group 502: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_Sample/req
      -- 
    req_3766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(502), ack => WPIPE_ConvTranspose_output_pipe_1454_inst_req_0); -- 
    convTranspose_cp_element_group_502: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_502"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(501) & convTranspose_CP_39_elements(467);
      gj_convTranspose_cp_element_group_502 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(502), clk => clk, reset => reset); --
    end block;
    -- CP-element group 503:  transition  input  output  bypass 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	502 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	504 
    -- CP-element group 503:  members (6) 
      -- CP-element group 503: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_sample_completed_
      -- CP-element group 503: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_update_start_
      -- CP-element group 503: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_Sample/$exit
      -- CP-element group 503: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_Sample/ack
      -- CP-element group 503: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_Update/req
      -- 
    ack_3767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 503_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0, ack => convTranspose_CP_39_elements(503)); -- 
    req_3771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(503), ack => WPIPE_ConvTranspose_output_pipe_1454_inst_req_1); -- 
    -- CP-element group 504:  transition  input  bypass 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	503 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	505 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_update_completed_
      -- CP-element group 504: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_Update/$exit
      -- CP-element group 504: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/WPIPE_ConvTranspose_output_pipe_1454_Update/ack
      -- 
    ack_3772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1, ack => convTranspose_CP_39_elements(504)); -- 
    -- CP-element group 505:  branch  join  transition  place  output  bypass 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	460 
    -- CP-element group 505: 	504 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	506 
    -- CP-element group 505: 	507 
    -- CP-element group 505:  members (10) 
      -- CP-element group 505: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467__exit__
      -- CP-element group 505: 	 branch_block_stmt_32/if_stmt_1468__entry__
      -- CP-element group 505: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/$exit
      -- CP-element group 505: 	 branch_block_stmt_32/if_stmt_1468_dead_link/$entry
      -- CP-element group 505: 	 branch_block_stmt_32/if_stmt_1468_eval_test/$entry
      -- CP-element group 505: 	 branch_block_stmt_32/if_stmt_1468_eval_test/$exit
      -- CP-element group 505: 	 branch_block_stmt_32/if_stmt_1468_eval_test/branch_req
      -- CP-element group 505: 	 branch_block_stmt_32/R_exitcond1_1469_place
      -- CP-element group 505: 	 branch_block_stmt_32/if_stmt_1468_if_link/$entry
      -- CP-element group 505: 	 branch_block_stmt_32/if_stmt_1468_else_link/$entry
      -- 
    branch_req_3780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(505), ack => if_stmt_1468_branch_req_0); -- 
    convTranspose_cp_element_group_505: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_505"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(460) & convTranspose_CP_39_elements(504);
      gj_convTranspose_cp_element_group_505 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(505), clk => clk, reset => reset); --
    end block;
    -- CP-element group 506:  merge  transition  place  input  bypass 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	505 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	535 
    -- CP-element group 506:  members (13) 
      -- CP-element group 506: 	 branch_block_stmt_32/merge_stmt_1474__exit__
      -- CP-element group 506: 	 branch_block_stmt_32/forx_xend702x_xloopexit_forx_xend702
      -- CP-element group 506: 	 branch_block_stmt_32/merge_stmt_1474_PhiAck/$exit
      -- CP-element group 506: 	 branch_block_stmt_32/forx_xend702x_xloopexit_forx_xend702_PhiReq/$entry
      -- CP-element group 506: 	 branch_block_stmt_32/forx_xend702x_xloopexit_forx_xend702_PhiReq/$exit
      -- CP-element group 506: 	 branch_block_stmt_32/merge_stmt_1474_PhiAck/$entry
      -- CP-element group 506: 	 branch_block_stmt_32/merge_stmt_1474_PhiAck/dummy
      -- CP-element group 506: 	 branch_block_stmt_32/merge_stmt_1474_PhiReqMerge
      -- CP-element group 506: 	 branch_block_stmt_32/forx_xbody630_forx_xend702x_xloopexit_PhiReq/$exit
      -- CP-element group 506: 	 branch_block_stmt_32/forx_xbody630_forx_xend702x_xloopexit_PhiReq/$entry
      -- CP-element group 506: 	 branch_block_stmt_32/if_stmt_1468_if_link/$exit
      -- CP-element group 506: 	 branch_block_stmt_32/if_stmt_1468_if_link/if_choice_transition
      -- CP-element group 506: 	 branch_block_stmt_32/forx_xbody630_forx_xend702x_xloopexit
      -- 
    if_choice_transition_3785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1468_branch_ack_1, ack => convTranspose_CP_39_elements(506)); -- 
    -- CP-element group 507:  fork  transition  place  input  output  bypass 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	505 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	530 
    -- CP-element group 507: 	531 
    -- CP-element group 507:  members (12) 
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/$entry
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/$entry
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/$entry
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/$entry
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/Update/cr
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/Sample/rr
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/$entry
      -- CP-element group 507: 	 branch_block_stmt_32/if_stmt_1468_else_link/$exit
      -- CP-element group 507: 	 branch_block_stmt_32/if_stmt_1468_else_link/else_choice_transition
      -- CP-element group 507: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630
      -- 
    else_choice_transition_3789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 507_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1468_branch_ack_0, ack => convTranspose_CP_39_elements(507)); -- 
    cr_4069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(507), ack => type_cast_1346_inst_req_1); -- 
    rr_4064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(507), ack => type_cast_1346_inst_req_0); -- 
    -- CP-element group 508:  merge  branch  transition  place  output  bypass 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	91 
    -- CP-element group 508: 	136 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	92 
    -- CP-element group 508: 	93 
    -- CP-element group 508:  members (17) 
      -- CP-element group 508: 	 branch_block_stmt_32/merge_stmt_358__exit__
      -- CP-element group 508: 	 branch_block_stmt_32/assign_stmt_364__entry__
      -- CP-element group 508: 	 branch_block_stmt_32/assign_stmt_364__exit__
      -- CP-element group 508: 	 branch_block_stmt_32/if_stmt_365__entry__
      -- CP-element group 508: 	 branch_block_stmt_32/assign_stmt_364/$entry
      -- CP-element group 508: 	 branch_block_stmt_32/assign_stmt_364/$exit
      -- CP-element group 508: 	 branch_block_stmt_32/if_stmt_365_dead_link/$entry
      -- CP-element group 508: 	 branch_block_stmt_32/if_stmt_365_eval_test/$entry
      -- CP-element group 508: 	 branch_block_stmt_32/if_stmt_365_eval_test/$exit
      -- CP-element group 508: 	 branch_block_stmt_32/if_stmt_365_eval_test/branch_req
      -- CP-element group 508: 	 branch_block_stmt_32/R_cmp194759_366_place
      -- CP-element group 508: 	 branch_block_stmt_32/if_stmt_365_if_link/$entry
      -- CP-element group 508: 	 branch_block_stmt_32/if_stmt_365_else_link/$entry
      -- CP-element group 508: 	 branch_block_stmt_32/merge_stmt_358_PhiReqMerge
      -- CP-element group 508: 	 branch_block_stmt_32/merge_stmt_358_PhiAck/$entry
      -- CP-element group 508: 	 branch_block_stmt_32/merge_stmt_358_PhiAck/$exit
      -- CP-element group 508: 	 branch_block_stmt_32/merge_stmt_358_PhiAck/dummy
      -- 
    branch_req_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(508), ack => if_stmt_365_branch_req_0); -- 
    convTranspose_CP_39_elements(508) <= OrReduce(convTranspose_CP_39_elements(91) & convTranspose_CP_39_elements(136));
    -- CP-element group 509:  transition  output  delay-element  bypass 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	95 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	513 
    -- CP-element group 509:  members (5) 
      -- CP-element group 509: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody_PhiReq/$exit
      -- CP-element group 509: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody_PhiReq/phi_stmt_403/$exit
      -- CP-element group 509: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/$exit
      -- CP-element group 509: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_407_konst_delay_trans
      -- CP-element group 509: 	 branch_block_stmt_32/bbx_xnph765_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_req
      -- 
    phi_stmt_403_req_3837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_403_req_3837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(509), ack => phi_stmt_403_req_0); -- 
    -- Element group convTranspose_CP_39_elements(509) is a control-delay.
    cp_element_509_delay: control_delay_element  generic map(name => " 509_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(95), ack => convTranspose_CP_39_elements(509), clk => clk, reset =>reset);
    -- CP-element group 510:  transition  input  bypass 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	137 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	512 
    -- CP-element group 510:  members (2) 
      -- CP-element group 510: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/Sample/$exit
      -- CP-element group 510: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/Sample/ra
      -- 
    ra_3857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 510_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_409_inst_ack_0, ack => convTranspose_CP_39_elements(510)); -- 
    -- CP-element group 511:  transition  input  bypass 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	137 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	512 
    -- CP-element group 511:  members (2) 
      -- CP-element group 511: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/Update/$exit
      -- CP-element group 511: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/Update/ca
      -- 
    ca_3862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 511_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_409_inst_ack_1, ack => convTranspose_CP_39_elements(511)); -- 
    -- CP-element group 512:  join  transition  output  bypass 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	510 
    -- CP-element group 512: 	511 
    -- CP-element group 512: successors 
    -- CP-element group 512: 	513 
    -- CP-element group 512:  members (6) 
      -- CP-element group 512: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 512: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/$exit
      -- CP-element group 512: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/$exit
      -- CP-element group 512: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/$exit
      -- CP-element group 512: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_sources/type_cast_409/SplitProtocol/$exit
      -- CP-element group 512: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_403/phi_stmt_403_req
      -- 
    phi_stmt_403_req_3863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_403_req_3863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(512), ack => phi_stmt_403_req_1); -- 
    convTranspose_cp_element_group_512: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_512"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(510) & convTranspose_CP_39_elements(511);
      gj_convTranspose_cp_element_group_512 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(512), clk => clk, reset => reset); --
    end block;
    -- CP-element group 513:  merge  transition  place  bypass 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	509 
    -- CP-element group 513: 	512 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	514 
    -- CP-element group 513:  members (2) 
      -- CP-element group 513: 	 branch_block_stmt_32/merge_stmt_402_PhiReqMerge
      -- CP-element group 513: 	 branch_block_stmt_32/merge_stmt_402_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(513) <= OrReduce(convTranspose_CP_39_elements(509) & convTranspose_CP_39_elements(512));
    -- CP-element group 514:  fork  transition  place  input  output  bypass 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	513 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	96 
    -- CP-element group 514: 	97 
    -- CP-element group 514: 	99 
    -- CP-element group 514: 	100 
    -- CP-element group 514: 	103 
    -- CP-element group 514: 	107 
    -- CP-element group 514: 	111 
    -- CP-element group 514: 	115 
    -- CP-element group 514: 	119 
    -- CP-element group 514: 	123 
    -- CP-element group 514: 	127 
    -- CP-element group 514: 	131 
    -- CP-element group 514: 	134 
    -- CP-element group 514:  members (56) 
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_32/merge_stmt_402__exit__
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565__entry__
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_526_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Update/word_access_complete/word_0/cr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Update/word_access_complete/word_0/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Update/word_access_complete/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/ptr_deref_552_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_508_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_resized_1
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_scaled_1
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_computed_1
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_resize_1/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_resize_1/$exit
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_resize_1/index_resize_req
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_resize_1/index_resize_ack
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_scale_1/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_scale_1/$exit
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_scale_1/scale_rename_req
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_index_scale_1/scale_rename_ack
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_update_start
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_Sample/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_Sample/req
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/array_obj_ref_415_final_index_sum_regn_Update/req
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_complete/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/addr_of_416_complete/req
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_sample_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_Sample/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/RPIPE_ConvTranspose_input_pipe_419_Sample/rr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_544_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_423_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_490_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_436_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_Update/$entry
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_454_Update/cr
      -- CP-element group 514: 	 branch_block_stmt_32/assign_stmt_417_to_assign_stmt_565/type_cast_472_update_start_
      -- CP-element group 514: 	 branch_block_stmt_32/merge_stmt_402_PhiAck/$exit
      -- CP-element group 514: 	 branch_block_stmt_32/merge_stmt_402_PhiAck/phi_stmt_403_ack
      -- 
    phi_stmt_403_ack_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 514_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_403_ack_0, ack => convTranspose_CP_39_elements(514)); -- 
    cr_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_472_inst_req_1); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_526_inst_req_1); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_508_inst_req_1); -- 
    cr_1121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => ptr_deref_552_store_0_req_1); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_544_inst_req_1); -- 
    req_827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => array_obj_ref_415_index_offset_req_0); -- 
    req_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => array_obj_ref_415_index_offset_req_1); -- 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => addr_of_416_final_reg_req_1); -- 
    rr_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => RPIPE_ConvTranspose_input_pipe_419_inst_req_0); -- 
    cr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_423_inst_req_1); -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_490_inst_req_1); -- 
    cr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_436_inst_req_1); -- 
    cr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(514), ack => type_cast_454_inst_req_1); -- 
    -- CP-element group 515:  transition  output  delay-element  bypass 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	139 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	519 
    -- CP-element group 515:  members (5) 
      -- CP-element group 515: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196_PhiReq/$exit
      -- CP-element group 515: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196_PhiReq/phi_stmt_610/$exit
      -- CP-element group 515: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/$exit
      -- CP-element group 515: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_614_konst_delay_trans
      -- CP-element group 515: 	 branch_block_stmt_32/bbx_xnph761_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_req
      -- 
    phi_stmt_610_req_3891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_610_req_3891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(515), ack => phi_stmt_610_req_0); -- 
    -- Element group convTranspose_CP_39_elements(515) is a control-delay.
    cp_element_515_delay: control_delay_element  generic map(name => " 515_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(139), ack => convTranspose_CP_39_elements(515), clk => clk, reset =>reset);
    -- CP-element group 516:  transition  input  bypass 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	181 
    -- CP-element group 516: successors 
    -- CP-element group 516: 	518 
    -- CP-element group 516:  members (2) 
      -- CP-element group 516: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/Sample/$exit
      -- CP-element group 516: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/Sample/ra
      -- 
    ra_3911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_0, ack => convTranspose_CP_39_elements(516)); -- 
    -- CP-element group 517:  transition  input  bypass 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	181 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	518 
    -- CP-element group 517:  members (2) 
      -- CP-element group 517: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/Update/$exit
      -- CP-element group 517: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/Update/ca
      -- 
    ca_3916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_1, ack => convTranspose_CP_39_elements(517)); -- 
    -- CP-element group 518:  join  transition  output  bypass 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	516 
    -- CP-element group 518: 	517 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	519 
    -- CP-element group 518:  members (6) 
      -- CP-element group 518: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 518: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/$exit
      -- CP-element group 518: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/$exit
      -- CP-element group 518: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/$exit
      -- CP-element group 518: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_sources/type_cast_616/SplitProtocol/$exit
      -- CP-element group 518: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_610/phi_stmt_610_req
      -- 
    phi_stmt_610_req_3917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_610_req_3917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(518), ack => phi_stmt_610_req_1); -- 
    convTranspose_cp_element_group_518: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_518"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(516) & convTranspose_CP_39_elements(517);
      gj_convTranspose_cp_element_group_518 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(518), clk => clk, reset => reset); --
    end block;
    -- CP-element group 519:  merge  transition  place  bypass 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	515 
    -- CP-element group 519: 	518 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	520 
    -- CP-element group 519:  members (2) 
      -- CP-element group 519: 	 branch_block_stmt_32/merge_stmt_609_PhiReqMerge
      -- CP-element group 519: 	 branch_block_stmt_32/merge_stmt_609_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(519) <= OrReduce(convTranspose_CP_39_elements(515) & convTranspose_CP_39_elements(518));
    -- CP-element group 520:  fork  transition  place  input  output  bypass 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	519 
    -- CP-element group 520: successors 
    -- CP-element group 520: 	175 
    -- CP-element group 520: 	178 
    -- CP-element group 520: 	171 
    -- CP-element group 520: 	155 
    -- CP-element group 520: 	159 
    -- CP-element group 520: 	163 
    -- CP-element group 520: 	167 
    -- CP-element group 520: 	151 
    -- CP-element group 520: 	140 
    -- CP-element group 520: 	141 
    -- CP-element group 520: 	143 
    -- CP-element group 520: 	144 
    -- CP-element group 520: 	147 
    -- CP-element group 520:  members (56) 
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/merge_stmt_609__exit__
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772__entry__
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_733_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_715_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_Update/req
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_Sample/req
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_Sample/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_final_index_sum_regn_update_start
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_Sample/rr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_679_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_Sample/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_scale_1/scale_rename_ack
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_scale_1/scale_rename_req
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_697_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_scale_1/$exit
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_scale_1/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_resize_1/index_resize_ack
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_resize_1/index_resize_req
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_resize_1/$exit
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_resize_1/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_computed_1
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_scaled_1
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/RPIPE_ConvTranspose_input_pipe_626_sample_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/array_obj_ref_622_index_resized_1
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_643_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_661_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_complete/req
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_630_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/addr_of_623_complete/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/type_cast_751_Update/cr
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_update_start_
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Update/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Update/word_access_complete/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Update/word_access_complete/word_0/$entry
      -- CP-element group 520: 	 branch_block_stmt_32/assign_stmt_624_to_assign_stmt_772/ptr_deref_759_Update/word_access_complete/word_0/cr
      -- CP-element group 520: 	 branch_block_stmt_32/merge_stmt_609_PhiAck/$exit
      -- CP-element group 520: 	 branch_block_stmt_32/merge_stmt_609_PhiAck/phi_stmt_610_ack
      -- 
    phi_stmt_610_ack_3922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_610_ack_0, ack => convTranspose_CP_39_elements(520)); -- 
    cr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => type_cast_733_inst_req_1); -- 
    cr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => type_cast_715_inst_req_1); -- 
    cr_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => type_cast_643_inst_req_1); -- 
    req_1191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => array_obj_ref_622_index_offset_req_1); -- 
    cr_1318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => type_cast_679_inst_req_1); -- 
    req_1186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => array_obj_ref_622_index_offset_req_0); -- 
    rr_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => RPIPE_ConvTranspose_input_pipe_626_inst_req_0); -- 
    cr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => type_cast_697_inst_req_1); -- 
    cr_1234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => type_cast_630_inst_req_1); -- 
    cr_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => type_cast_661_inst_req_1); -- 
    req_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => addr_of_623_final_reg_req_1); -- 
    cr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => type_cast_751_inst_req_1); -- 
    cr_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(520), ack => ptr_deref_759_store_0_req_1); -- 
    -- CP-element group 521:  merge  branch  transition  place  output  bypass 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	180 
    -- CP-element group 521: 	93 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	182 
    -- CP-element group 521: 	183 
    -- CP-element group 521:  members (17) 
      -- CP-element group 521: 	 branch_block_stmt_32/merge_stmt_781__exit__
      -- CP-element group 521: 	 branch_block_stmt_32/assign_stmt_786_to_assign_stmt_797__entry__
      -- CP-element group 521: 	 branch_block_stmt_32/assign_stmt_786_to_assign_stmt_797__exit__
      -- CP-element group 521: 	 branch_block_stmt_32/if_stmt_798__entry__
      -- CP-element group 521: 	 branch_block_stmt_32/assign_stmt_786_to_assign_stmt_797/$entry
      -- CP-element group 521: 	 branch_block_stmt_32/assign_stmt_786_to_assign_stmt_797/$exit
      -- CP-element group 521: 	 branch_block_stmt_32/if_stmt_798_dead_link/$entry
      -- CP-element group 521: 	 branch_block_stmt_32/if_stmt_798_eval_test/$entry
      -- CP-element group 521: 	 branch_block_stmt_32/if_stmt_798_eval_test/$exit
      -- CP-element group 521: 	 branch_block_stmt_32/if_stmt_798_eval_test/branch_req
      -- CP-element group 521: 	 branch_block_stmt_32/R_cmp264755_799_place
      -- CP-element group 521: 	 branch_block_stmt_32/if_stmt_798_if_link/$entry
      -- CP-element group 521: 	 branch_block_stmt_32/if_stmt_798_else_link/$entry
      -- CP-element group 521: 	 branch_block_stmt_32/merge_stmt_781_PhiReqMerge
      -- CP-element group 521: 	 branch_block_stmt_32/merge_stmt_781_PhiAck/$entry
      -- CP-element group 521: 	 branch_block_stmt_32/merge_stmt_781_PhiAck/$exit
      -- CP-element group 521: 	 branch_block_stmt_32/merge_stmt_781_PhiAck/dummy
      -- 
    branch_req_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(521), ack => if_stmt_798_branch_req_0); -- 
    convTranspose_CP_39_elements(521) <= OrReduce(convTranspose_CP_39_elements(180) & convTranspose_CP_39_elements(93));
    -- CP-element group 522:  transition  output  delay-element  bypass 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	185 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	526 
    -- CP-element group 522:  members (5) 
      -- CP-element group 522: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266_PhiReq/$exit
      -- CP-element group 522: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266_PhiReq/phi_stmt_842/$exit
      -- CP-element group 522: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/$exit
      -- CP-element group 522: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_846_konst_delay_trans
      -- CP-element group 522: 	 branch_block_stmt_32/bbx_xnph757_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_req
      -- 
    phi_stmt_842_req_3968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_842_req_3968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(522), ack => phi_stmt_842_req_0); -- 
    -- Element group convTranspose_CP_39_elements(522) is a control-delay.
    cp_element_522_delay: control_delay_element  generic map(name => " 522_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(185), ack => convTranspose_CP_39_elements(522), clk => clk, reset =>reset);
    -- CP-element group 523:  transition  input  bypass 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	194 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	525 
    -- CP-element group 523:  members (2) 
      -- CP-element group 523: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/Sample/$exit
      -- CP-element group 523: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/Sample/ra
      -- 
    ra_3988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 523_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_848_inst_ack_0, ack => convTranspose_CP_39_elements(523)); -- 
    -- CP-element group 524:  transition  input  bypass 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	194 
    -- CP-element group 524: successors 
    -- CP-element group 524: 	525 
    -- CP-element group 524:  members (2) 
      -- CP-element group 524: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/Update/$exit
      -- CP-element group 524: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/Update/ca
      -- 
    ca_3993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_848_inst_ack_1, ack => convTranspose_CP_39_elements(524)); -- 
    -- CP-element group 525:  join  transition  output  bypass 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	523 
    -- CP-element group 525: 	524 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	526 
    -- CP-element group 525:  members (6) 
      -- CP-element group 525: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 525: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/$exit
      -- CP-element group 525: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/$exit
      -- CP-element group 525: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/$exit
      -- CP-element group 525: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_sources/type_cast_848/SplitProtocol/$exit
      -- CP-element group 525: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_842/phi_stmt_842_req
      -- 
    phi_stmt_842_req_3994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_842_req_3994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(525), ack => phi_stmt_842_req_1); -- 
    convTranspose_cp_element_group_525: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_525"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(523) & convTranspose_CP_39_elements(524);
      gj_convTranspose_cp_element_group_525 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(525), clk => clk, reset => reset); --
    end block;
    -- CP-element group 526:  merge  transition  place  bypass 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	522 
    -- CP-element group 526: 	525 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	527 
    -- CP-element group 526:  members (2) 
      -- CP-element group 526: 	 branch_block_stmt_32/merge_stmt_841_PhiReqMerge
      -- CP-element group 526: 	 branch_block_stmt_32/merge_stmt_841_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(526) <= OrReduce(convTranspose_CP_39_elements(522) & convTranspose_CP_39_elements(525));
    -- CP-element group 527:  fork  transition  place  input  output  bypass 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	526 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	186 
    -- CP-element group 527: 	187 
    -- CP-element group 527: 	189 
    -- CP-element group 527: 	191 
    -- CP-element group 527:  members (29) 
      -- CP-element group 527: 	 branch_block_stmt_32/merge_stmt_841__exit__
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872__entry__
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_update_start_
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_resized_1
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_scaled_1
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_computed_1
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_resize_1/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_resize_1/$exit
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_resize_1/index_resize_req
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_resize_1/index_resize_ack
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_scale_1/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_scale_1/$exit
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_scale_1/scale_rename_req
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_index_scale_1/scale_rename_ack
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_update_start
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_Sample/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_Sample/req
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/array_obj_ref_854_final_index_sum_regn_Update/req
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_complete/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/addr_of_855_complete/req
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_update_start_
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Update/word_access_complete/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Update/word_access_complete/word_0/$entry
      -- CP-element group 527: 	 branch_block_stmt_32/assign_stmt_856_to_assign_stmt_872/ptr_deref_858_Update/word_access_complete/word_0/cr
      -- CP-element group 527: 	 branch_block_stmt_32/merge_stmt_841_PhiAck/$exit
      -- CP-element group 527: 	 branch_block_stmt_32/merge_stmt_841_PhiAck/phi_stmt_842_ack
      -- 
    phi_stmt_842_ack_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_842_ack_0, ack => convTranspose_CP_39_elements(527)); -- 
    req_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => array_obj_ref_854_index_offset_req_0); -- 
    req_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => array_obj_ref_854_index_offset_req_1); -- 
    req_1587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => addr_of_855_final_reg_req_1); -- 
    cr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(527), ack => ptr_deref_858_store_0_req_1); -- 
    -- CP-element group 528:  merge  fork  transition  place  output  bypass 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	183 
    -- CP-element group 528: 	193 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	195 
    -- CP-element group 528: 	196 
    -- CP-element group 528: 	198 
    -- CP-element group 528: 	199 
    -- CP-element group 528: 	255 
    -- CP-element group 528: 	291 
    -- CP-element group 528: 	292 
    -- CP-element group 528: 	296 
    -- CP-element group 528: 	297 
    -- CP-element group 528: 	319 
    -- CP-element group 528: 	357 
    -- CP-element group 528: 	358 
    -- CP-element group 528: 	380 
    -- CP-element group 528: 	418 
    -- CP-element group 528: 	419 
    -- CP-element group 528: 	441 
    -- CP-element group 528: 	443 
    -- CP-element group 528: 	445 
    -- CP-element group 528: 	447 
    -- CP-element group 528:  members (64) 
      -- CP-element group 528: 	 branch_block_stmt_32/merge_stmt_881__exit__
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278__entry__
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_Update/cr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_update_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_Sample/crr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/call_stmt_884_Update/ccr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_update_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_889_Update/cr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_update_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block0_start_891_Sample/req
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1035_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_Update/cr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_Sample/req
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_update_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1048_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block3_done_1277_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block1_start_979_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block2_start_1077_Sample/req
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_Update/cr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_update_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block2_done_1274_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1238_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_update_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block0_done_1268_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_Sample/rr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_Update/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/type_cast_1143_Update/cr
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/RPIPE_Block1_done_1271_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_sample_start_
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_Sample/$entry
      -- CP-element group 528: 	 branch_block_stmt_32/call_stmt_884_to_assign_stmt_1278/WPIPE_Block3_start_1172_Sample/req
      -- CP-element group 528: 	 branch_block_stmt_32/merge_stmt_881_PhiAck/dummy
      -- CP-element group 528: 	 branch_block_stmt_32/merge_stmt_881_PhiReqMerge
      -- CP-element group 528: 	 branch_block_stmt_32/merge_stmt_881_PhiAck/$exit
      -- CP-element group 528: 	 branch_block_stmt_32/merge_stmt_881_PhiAck/$entry
      -- 
    cr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_1035_inst_req_1); -- 
    rr_3320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => RPIPE_Block0_done_1268_inst_req_0); -- 
    rr_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_1035_inst_req_0); -- 
    crr_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => call_stmt_884_call_req_0); -- 
    ccr_1673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => call_stmt_884_call_req_1); -- 
    cr_1687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_889_inst_req_1); -- 
    req_1696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => WPIPE_Block0_start_891_inst_req_0); -- 
    cr_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_1048_inst_req_1); -- 
    rr_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_1048_inst_req_0); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => WPIPE_Block1_start_979_inst_req_0); -- 
    rr_3362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => RPIPE_Block3_done_1277_inst_req_0); -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => WPIPE_Block2_start_1077_inst_req_0); -- 
    cr_3185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_1238_inst_req_1); -- 
    rr_3348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => RPIPE_Block2_done_1274_inst_req_0); -- 
    rr_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_1238_inst_req_0); -- 
    rr_3334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => RPIPE_Block1_done_1271_inst_req_0); -- 
    rr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_1143_inst_req_0); -- 
    cr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => type_cast_1143_inst_req_1); -- 
    req_2914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(528), ack => WPIPE_Block3_start_1172_inst_req_0); -- 
    convTranspose_CP_39_elements(528) <= OrReduce(convTranspose_CP_39_elements(183) & convTranspose_CP_39_elements(193));
    -- CP-element group 529:  transition  output  delay-element  bypass 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	459 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	533 
    -- CP-element group 529:  members (5) 
      -- CP-element group 529: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630_PhiReq/$exit
      -- CP-element group 529: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_req
      -- CP-element group 529: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1344_konst_delay_trans
      -- CP-element group 529: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/$exit
      -- CP-element group 529: 	 branch_block_stmt_32/bbx_xnph_forx_xbody630_PhiReq/phi_stmt_1340/$exit
      -- 
    phi_stmt_1340_req_4045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1340_req_4045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(529), ack => phi_stmt_1340_req_0); -- 
    -- Element group convTranspose_CP_39_elements(529) is a control-delay.
    cp_element_529_delay: control_delay_element  generic map(name => " 529_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(459), ack => convTranspose_CP_39_elements(529), clk => clk, reset =>reset);
    -- CP-element group 530:  transition  input  bypass 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	507 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	532 
    -- CP-element group 530:  members (2) 
      -- CP-element group 530: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/Sample/ra
      -- CP-element group 530: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/Sample/$exit
      -- 
    ra_4065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 530_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_0, ack => convTranspose_CP_39_elements(530)); -- 
    -- CP-element group 531:  transition  input  bypass 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	507 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	532 
    -- CP-element group 531:  members (2) 
      -- CP-element group 531: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/Update/ca
      -- CP-element group 531: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/Update/$exit
      -- 
    ca_4070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1346_inst_ack_1, ack => convTranspose_CP_39_elements(531)); -- 
    -- CP-element group 532:  join  transition  output  bypass 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	530 
    -- CP-element group 532: 	531 
    -- CP-element group 532: successors 
    -- CP-element group 532: 	533 
    -- CP-element group 532:  members (6) 
      -- CP-element group 532: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/$exit
      -- CP-element group 532: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/$exit
      -- CP-element group 532: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/$exit
      -- CP-element group 532: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/$exit
      -- CP-element group 532: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_req
      -- CP-element group 532: 	 branch_block_stmt_32/forx_xbody630_forx_xbody630_PhiReq/phi_stmt_1340/phi_stmt_1340_sources/type_cast_1346/SplitProtocol/$exit
      -- 
    phi_stmt_1340_req_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1340_req_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(532), ack => phi_stmt_1340_req_1); -- 
    convTranspose_cp_element_group_532: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_532"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(530) & convTranspose_CP_39_elements(531);
      gj_convTranspose_cp_element_group_532 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(532), clk => clk, reset => reset); --
    end block;
    -- CP-element group 533:  merge  transition  place  bypass 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	529 
    -- CP-element group 533: 	532 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	534 
    -- CP-element group 533:  members (2) 
      -- CP-element group 533: 	 branch_block_stmt_32/merge_stmt_1339_PhiReqMerge
      -- CP-element group 533: 	 branch_block_stmt_32/merge_stmt_1339_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(533) <= OrReduce(convTranspose_CP_39_elements(529) & convTranspose_CP_39_elements(532));
    -- CP-element group 534:  fork  transition  place  input  output  bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	533 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	460 
    -- CP-element group 534: 	461 
    -- CP-element group 534: 	463 
    -- CP-element group 534: 	471 
    -- CP-element group 534: 	473 
    -- CP-element group 534: 	475 
    -- CP-element group 534: 	477 
    -- CP-element group 534: 	479 
    -- CP-element group 534: 	481 
    -- CP-element group 534: 	465 
    -- CP-element group 534: 	467 
    -- CP-element group 534: 	469 
    -- CP-element group 534:  members (53) 
      -- CP-element group 534: 	 branch_block_stmt_32/merge_stmt_1339__exit__
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467__entry__
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_resized_1
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_scaled_1
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_computed_1
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_resize_1/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_resize_1/$exit
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_resize_1/index_resize_req
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_resize_1/index_resize_ack
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_scale_1/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_scale_1/$exit
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_scale_1/scale_rename_req
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_index_scale_1/scale_rename_ack
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_update_start
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_Sample/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_Sample/req
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/array_obj_ref_1352_final_index_sum_regn_Update/req
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_complete/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/addr_of_1353_complete/req
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/word_access_complete/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/word_access_complete/word_0/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/ptr_deref_1357_Update/word_access_complete/word_0/cr
      -- CP-element group 534: 	 branch_block_stmt_32/merge_stmt_1339_PhiAck/phi_stmt_1340_ack
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1361_Update/cr
      -- CP-element group 534: 	 branch_block_stmt_32/merge_stmt_1339_PhiAck/$exit
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1371_Update/cr
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1381_Update/cr
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1391_Update/cr
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1401_Update/cr
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1411_Update/cr
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1421_Update/cr
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_update_start_
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_32/assign_stmt_1354_to_assign_stmt_1467/type_cast_1431_Update/cr
      -- 
    phi_stmt_1340_ack_4076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1340_ack_0, ack => convTranspose_CP_39_elements(534)); -- 
    req_3477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => array_obj_ref_1352_index_offset_req_0); -- 
    req_3482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => array_obj_ref_1352_index_offset_req_1); -- 
    req_3497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => addr_of_1353_final_reg_req_1); -- 
    cr_3542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => ptr_deref_1357_load_0_req_1); -- 
    cr_3561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => type_cast_1361_inst_req_1); -- 
    cr_3575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => type_cast_1371_inst_req_1); -- 
    cr_3589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => type_cast_1381_inst_req_1); -- 
    cr_3603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => type_cast_1391_inst_req_1); -- 
    cr_3617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => type_cast_1401_inst_req_1); -- 
    cr_3631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => type_cast_1411_inst_req_1); -- 
    cr_3645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => type_cast_1421_inst_req_1); -- 
    cr_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(534), ack => type_cast_1431_inst_req_1); -- 
    -- CP-element group 535:  merge  transition  place  bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	506 
    -- CP-element group 535: 	457 
    -- CP-element group 535: successors 
    -- CP-element group 535:  members (16) 
      -- CP-element group 535: 	 $exit
      -- CP-element group 535: 	 branch_block_stmt_32/$exit
      -- CP-element group 535: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1476__exit__
      -- CP-element group 535: 	 branch_block_stmt_32/return__
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1478__exit__
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1476_PhiReqMerge
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1478_PhiReqMerge
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1476_PhiAck/$entry
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1476_PhiAck/$exit
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1476_PhiAck/dummy
      -- CP-element group 535: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 535: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1478_PhiAck/$entry
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1478_PhiAck/$exit
      -- CP-element group 535: 	 branch_block_stmt_32/merge_stmt_1478_PhiAck/dummy
      -- 
    convTranspose_CP_39_elements(535) <= OrReduce(convTranspose_CP_39_elements(506) & convTranspose_CP_39_elements(457));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar772_853_resized : std_logic_vector(13 downto 0);
    signal R_indvar772_853_scaled : std_logic_vector(13 downto 0);
    signal R_indvar783_621_resized : std_logic_vector(10 downto 0);
    signal R_indvar783_621_scaled : std_logic_vector(10 downto 0);
    signal R_indvar795_414_resized : std_logic_vector(13 downto 0);
    signal R_indvar795_414_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1351_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1351_scaled : std_logic_vector(13 downto 0);
    signal add117_292 : std_logic_vector(31 downto 0);
    signal add126_317 : std_logic_vector(31 downto 0);
    signal add12_82 : std_logic_vector(31 downto 0);
    signal add135_342 : std_logic_vector(31 downto 0);
    signal add150_442 : std_logic_vector(63 downto 0);
    signal add156_460 : std_logic_vector(63 downto 0);
    signal add162_478 : std_logic_vector(63 downto 0);
    signal add168_496 : std_logic_vector(63 downto 0);
    signal add174_514 : std_logic_vector(63 downto 0);
    signal add180_532 : std_logic_vector(63 downto 0);
    signal add186_550 : std_logic_vector(63 downto 0);
    signal add206_649 : std_logic_vector(63 downto 0);
    signal add212_667 : std_logic_vector(63 downto 0);
    signal add218_685 : std_logic_vector(63 downto 0);
    signal add21_107 : std_logic_vector(31 downto 0);
    signal add224_703 : std_logic_vector(63 downto 0);
    signal add230_721 : std_logic_vector(63 downto 0);
    signal add236_739 : std_logic_vector(63 downto 0);
    signal add242_757 : std_logic_vector(63 downto 0);
    signal add30_132 : std_logic_vector(31 downto 0);
    signal add39_157 : std_logic_vector(31 downto 0);
    signal add48_182 : std_logic_vector(31 downto 0);
    signal add57_207 : std_logic_vector(31 downto 0);
    signal add74_235 : std_logic_vector(31 downto 0);
    signal add79_240 : std_logic_vector(31 downto 0);
    signal add_57 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1352_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1352_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1352_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1352_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1352_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1352_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_415_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_622_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_622_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_622_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_622_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_622_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_622_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_854_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_854_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_854_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_854_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_854_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_854_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_624 : std_logic_vector(31 downto 0);
    signal arrayidx269_856 : std_logic_vector(31 downto 0);
    signal arrayidx635_1354 : std_logic_vector(31 downto 0);
    signal arrayidx_417 : std_logic_vector(31 downto 0);
    signal call101_264 : std_logic_vector(7 downto 0);
    signal call106_267 : std_logic_vector(7 downto 0);
    signal call10_73 : std_logic_vector(7 downto 0);
    signal call110_270 : std_logic_vector(7 downto 0);
    signal call115_283 : std_logic_vector(7 downto 0);
    signal call119_295 : std_logic_vector(7 downto 0);
    signal call124_308 : std_logic_vector(7 downto 0);
    signal call128_320 : std_logic_vector(7 downto 0);
    signal call133_333 : std_logic_vector(7 downto 0);
    signal call143_420 : std_logic_vector(7 downto 0);
    signal call147_433 : std_logic_vector(7 downto 0);
    signal call14_85 : std_logic_vector(7 downto 0);
    signal call153_451 : std_logic_vector(7 downto 0);
    signal call159_469 : std_logic_vector(7 downto 0);
    signal call165_487 : std_logic_vector(7 downto 0);
    signal call171_505 : std_logic_vector(7 downto 0);
    signal call177_523 : std_logic_vector(7 downto 0);
    signal call183_541 : std_logic_vector(7 downto 0);
    signal call199_627 : std_logic_vector(7 downto 0);
    signal call19_98 : std_logic_vector(7 downto 0);
    signal call203_640 : std_logic_vector(7 downto 0);
    signal call209_658 : std_logic_vector(7 downto 0);
    signal call215_676 : std_logic_vector(7 downto 0);
    signal call221_694 : std_logic_vector(7 downto 0);
    signal call227_712 : std_logic_vector(7 downto 0);
    signal call233_730 : std_logic_vector(7 downto 0);
    signal call239_748 : std_logic_vector(7 downto 0);
    signal call23_110 : std_logic_vector(7 downto 0);
    signal call275_884 : std_logic_vector(63 downto 0);
    signal call28_123 : std_logic_vector(7 downto 0);
    signal call2_48 : std_logic_vector(7 downto 0);
    signal call32_135 : std_logic_vector(7 downto 0);
    signal call37_148 : std_logic_vector(7 downto 0);
    signal call41_160 : std_logic_vector(7 downto 0);
    signal call46_173 : std_logic_vector(7 downto 0);
    signal call50_185 : std_logic_vector(7 downto 0);
    signal call55_198 : std_logic_vector(7 downto 0);
    signal call5_60 : std_logic_vector(7 downto 0);
    signal call610_1269 : std_logic_vector(7 downto 0);
    signal call612_1272 : std_logic_vector(7 downto 0);
    signal call614_1275 : std_logic_vector(7 downto 0);
    signal call616_1278 : std_logic_vector(7 downto 0);
    signal call618_1281 : std_logic_vector(63 downto 0);
    signal call92_258 : std_logic_vector(7 downto 0);
    signal call97_261 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp194759_364 : std_logic_vector(0 downto 0);
    signal cmp264755_797 : std_logic_vector(0 downto 0);
    signal cmp763_349 : std_logic_vector(0 downto 0);
    signal conv113_274 : std_logic_vector(31 downto 0);
    signal conv116_287 : std_logic_vector(31 downto 0);
    signal conv11_77 : std_logic_vector(31 downto 0);
    signal conv122_299 : std_logic_vector(31 downto 0);
    signal conv125_312 : std_logic_vector(31 downto 0);
    signal conv131_324 : std_logic_vector(31 downto 0);
    signal conv134_337 : std_logic_vector(31 downto 0);
    signal conv144_424 : std_logic_vector(63 downto 0);
    signal conv149_437 : std_logic_vector(63 downto 0);
    signal conv155_455 : std_logic_vector(63 downto 0);
    signal conv161_473 : std_logic_vector(63 downto 0);
    signal conv167_491 : std_logic_vector(63 downto 0);
    signal conv173_509 : std_logic_vector(63 downto 0);
    signal conv179_527 : std_logic_vector(63 downto 0);
    signal conv17_89 : std_logic_vector(31 downto 0);
    signal conv185_545 : std_logic_vector(63 downto 0);
    signal conv1_39 : std_logic_vector(31 downto 0);
    signal conv200_631 : std_logic_vector(63 downto 0);
    signal conv205_644 : std_logic_vector(63 downto 0);
    signal conv20_102 : std_logic_vector(31 downto 0);
    signal conv211_662 : std_logic_vector(63 downto 0);
    signal conv217_680 : std_logic_vector(63 downto 0);
    signal conv223_698 : std_logic_vector(63 downto 0);
    signal conv229_716 : std_logic_vector(63 downto 0);
    signal conv235_734 : std_logic_vector(63 downto 0);
    signal conv241_752 : std_logic_vector(63 downto 0);
    signal conv26_114 : std_logic_vector(31 downto 0);
    signal conv276_890 : std_logic_vector(63 downto 0);
    signal conv29_127 : std_logic_vector(31 downto 0);
    signal conv35_139 : std_logic_vector(31 downto 0);
    signal conv38_152 : std_logic_vector(31 downto 0);
    signal conv3_52 : std_logic_vector(31 downto 0);
    signal conv415_1036 : std_logic_vector(7 downto 0);
    signal conv418_1049 : std_logic_vector(7 downto 0);
    signal conv44_164 : std_logic_vector(31 downto 0);
    signal conv47_177 : std_logic_vector(31 downto 0);
    signal conv501_1144 : std_logic_vector(7 downto 0);
    signal conv53_189 : std_logic_vector(31 downto 0);
    signal conv56_202 : std_logic_vector(31 downto 0);
    signal conv584_1239 : std_logic_vector(7 downto 0);
    signal conv619_1286 : std_logic_vector(63 downto 0);
    signal conv639_1362 : std_logic_vector(7 downto 0);
    signal conv645_1372 : std_logic_vector(7 downto 0);
    signal conv651_1382 : std_logic_vector(7 downto 0);
    signal conv657_1392 : std_logic_vector(7 downto 0);
    signal conv663_1402 : std_logic_vector(7 downto 0);
    signal conv669_1412 : std_logic_vector(7 downto 0);
    signal conv675_1422 : std_logic_vector(7 downto 0);
    signal conv681_1432 : std_logic_vector(7 downto 0);
    signal conv8_64 : std_logic_vector(31 downto 0);
    signal exitcond1_1467 : std_logic_vector(0 downto 0);
    signal exitcond2_772 : std_logic_vector(0 downto 0);
    signal exitcond3_565 : std_logic_vector(0 downto 0);
    signal exitcond_872 : std_logic_vector(0 downto 0);
    signal iNsTr_14_229 : std_logic_vector(31 downto 0);
    signal iNsTr_26_387 : std_logic_vector(63 downto 0);
    signal iNsTr_292_1324 : std_logic_vector(63 downto 0);
    signal iNsTr_39_594 : std_logic_vector(63 downto 0);
    signal iNsTr_53_826 : std_logic_vector(63 downto 0);
    signal indvar772_842 : std_logic_vector(63 downto 0);
    signal indvar783_610 : std_logic_vector(63 downto 0);
    signal indvar795_403 : std_logic_vector(63 downto 0);
    signal indvar_1340 : std_logic_vector(63 downto 0);
    signal indvarx_xnext773_867 : std_logic_vector(63 downto 0);
    signal indvarx_xnext784_767 : std_logic_vector(63 downto 0);
    signal indvarx_xnext796_560 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1462 : std_logic_vector(63 downto 0);
    signal mul256_786 : std_logic_vector(31 downto 0);
    signal mul259_791 : std_logic_vector(31 downto 0);
    signal mul66_217 : std_logic_vector(31 downto 0);
    signal mul85_245 : std_logic_vector(31 downto 0);
    signal mul88_250 : std_logic_vector(31 downto 0);
    signal mul91_255 : std_logic_vector(31 downto 0);
    signal mul_212 : std_logic_vector(31 downto 0);
    signal ptr_deref_1357_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1357_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1357_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1357_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1357_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_552_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_552_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_552_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_552_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_552_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_552_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_759_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_759_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_759_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_759_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_759_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_759_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_858_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_858_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_858_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_858_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_858_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_858_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl114_280 : std_logic_vector(31 downto 0);
    signal shl123_305 : std_logic_vector(31 downto 0);
    signal shl132_330 : std_logic_vector(31 downto 0);
    signal shl146_430 : std_logic_vector(63 downto 0);
    signal shl152_448 : std_logic_vector(63 downto 0);
    signal shl158_466 : std_logic_vector(63 downto 0);
    signal shl164_484 : std_logic_vector(63 downto 0);
    signal shl170_502 : std_logic_vector(63 downto 0);
    signal shl176_520 : std_logic_vector(63 downto 0);
    signal shl182_538 : std_logic_vector(63 downto 0);
    signal shl18_95 : std_logic_vector(31 downto 0);
    signal shl202_637 : std_logic_vector(63 downto 0);
    signal shl208_655 : std_logic_vector(63 downto 0);
    signal shl214_673 : std_logic_vector(63 downto 0);
    signal shl220_691 : std_logic_vector(63 downto 0);
    signal shl226_709 : std_logic_vector(63 downto 0);
    signal shl232_727 : std_logic_vector(63 downto 0);
    signal shl238_745 : std_logic_vector(63 downto 0);
    signal shl27_120 : std_logic_vector(31 downto 0);
    signal shl36_145 : std_logic_vector(31 downto 0);
    signal shl45_170 : std_logic_vector(31 downto 0);
    signal shl54_195 : std_logic_vector(31 downto 0);
    signal shl9_70 : std_logic_vector(31 downto 0);
    signal shl_45 : std_logic_vector(31 downto 0);
    signal shr417_1045 : std_logic_vector(31 downto 0);
    signal shr500_1140 : std_logic_vector(31 downto 0);
    signal shr583_1235 : std_logic_vector(31 downto 0);
    signal shr642_1368 : std_logic_vector(63 downto 0);
    signal shr648_1378 : std_logic_vector(63 downto 0);
    signal shr654_1388 : std_logic_vector(63 downto 0);
    signal shr660_1398 : std_logic_vector(63 downto 0);
    signal shr666_1408 : std_logic_vector(63 downto 0);
    signal shr672_1418 : std_logic_vector(63 downto 0);
    signal shr678_1428 : std_logic_vector(63 downto 0);
    signal shr_223 : std_logic_vector(31 downto 0);
    signal sub_1291 : std_logic_vector(63 downto 0);
    signal tmp636_1358 : std_logic_vector(63 downto 0);
    signal tmp767_1308 : std_logic_vector(31 downto 0);
    signal tmp767x_xop_1320 : std_logic_vector(31 downto 0);
    signal tmp768_1314 : std_logic_vector(0 downto 0);
    signal tmp771_1337 : std_logic_vector(63 downto 0);
    signal tmp776_810 : std_logic_vector(31 downto 0);
    signal tmp776x_xop_822 : std_logic_vector(31 downto 0);
    signal tmp777_816 : std_logic_vector(0 downto 0);
    signal tmp781_839 : std_logic_vector(63 downto 0);
    signal tmp788_578 : std_logic_vector(31 downto 0);
    signal tmp788x_xop_590 : std_logic_vector(31 downto 0);
    signal tmp789_584 : std_logic_vector(0 downto 0);
    signal tmp793_607 : std_logic_vector(63 downto 0);
    signal tmp799x_xop_383 : std_logic_vector(31 downto 0);
    signal tmp800_377 : std_logic_vector(0 downto 0);
    signal tmp804_400 : std_logic_vector(63 downto 0);
    signal type_cast_1043_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1133_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1138_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1228_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1284_wire : std_logic_vector(63 downto 0);
    signal type_cast_1306_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1312_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1318_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1328_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1335_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1344_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1346_wire : std_logic_vector(63 downto 0);
    signal type_cast_1366_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1376_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1386_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1396_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1406_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1416_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1426_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_143_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1460_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_168_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_193_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_221_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_227_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_278_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_303_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_328_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_346_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_362_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_375_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_381_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_391_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_398_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_407_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_409_wire : std_logic_vector(63 downto 0);
    signal type_cast_428_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_43_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_446_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_464_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_482_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_500_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_518_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_536_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_558_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_576_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_588_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_598_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_605_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_614_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_616_wire : std_logic_vector(63 downto 0);
    signal type_cast_635_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_653_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_671_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_689_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_707_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_725_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_743_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_765_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_795_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_808_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_814_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_820_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_830_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_837_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_846_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_848_wire : std_logic_vector(63 downto 0);
    signal type_cast_860_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_865_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_888_wire : std_logic_vector(63 downto 0);
    signal type_cast_93_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_947_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_951_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_955_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_959_wire_constant : std_logic_vector(7 downto 0);
    signal xx_xop806_832 : std_logic_vector(63 downto 0);
    signal xx_xop807_600 : std_logic_vector(63 downto 0);
    signal xx_xop808_393 : std_logic_vector(63 downto 0);
    signal xx_xop_1330 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1352_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1352_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1352_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1352_resized_base_address <= "00000000000000";
    array_obj_ref_415_constant_part_of_offset <= "00000000000000";
    array_obj_ref_415_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_415_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_415_resized_base_address <= "00000000000000";
    array_obj_ref_622_constant_part_of_offset <= "00000100010";
    array_obj_ref_622_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_622_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_622_resized_base_address <= "00000000000";
    array_obj_ref_854_constant_part_of_offset <= "00000000000000";
    array_obj_ref_854_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_854_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_854_resized_base_address <= "00000000000000";
    ptr_deref_1357_word_offset_0 <= "00000000000000";
    ptr_deref_552_word_offset_0 <= "00000000000000";
    ptr_deref_759_word_offset_0 <= "00000000000";
    ptr_deref_858_word_offset_0 <= "00000000000000";
    type_cast_1043_wire_constant <= "00000000000000000000000000001010";
    type_cast_1133_wire_constant <= "00000000";
    type_cast_1138_wire_constant <= "00000000000000000000000000001001";
    type_cast_118_wire_constant <= "00000000000000000000000000001000";
    type_cast_1228_wire_constant <= "00000000";
    type_cast_1233_wire_constant <= "00000000000000000000000000001000";
    type_cast_1306_wire_constant <= "00000000000000000000000000000010";
    type_cast_1312_wire_constant <= "00000000000000000000000000000001";
    type_cast_1318_wire_constant <= "11111111111111111111111111111111";
    type_cast_1328_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1335_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1344_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1366_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1376_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1396_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1406_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1416_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1426_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_143_wire_constant <= "00000000000000000000000000001000";
    type_cast_1460_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_168_wire_constant <= "00000000000000000000000000001000";
    type_cast_193_wire_constant <= "00000000000000000000000000001000";
    type_cast_221_wire_constant <= "00000000000000000000000000000010";
    type_cast_227_wire_constant <= "00000000000000000000000000000001";
    type_cast_233_wire_constant <= "00000000000000001111111111111110";
    type_cast_278_wire_constant <= "00000000000000000000000000001000";
    type_cast_303_wire_constant <= "00000000000000000000000000001000";
    type_cast_328_wire_constant <= "00000000000000000000000000001000";
    type_cast_346_wire_constant <= "00000000000000000000000000000011";
    type_cast_362_wire_constant <= "00000000000000000000000000000011";
    type_cast_375_wire_constant <= "00000000000000000000000000000001";
    type_cast_381_wire_constant <= "11111111111111111111111111111111";
    type_cast_391_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_398_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_407_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_428_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_43_wire_constant <= "00000000000000000000000000001000";
    type_cast_446_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_464_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_482_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_500_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_518_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_536_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_558_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_576_wire_constant <= "00000000000000000000000000000010";
    type_cast_582_wire_constant <= "00000000000000000000000000000001";
    type_cast_588_wire_constant <= "11111111111111111111111111111111";
    type_cast_598_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_605_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_614_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_635_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_653_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_671_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_689_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_68_wire_constant <= "00000000000000000000000000001000";
    type_cast_707_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_725_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_743_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_765_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_795_wire_constant <= "00000000000000000000000000000011";
    type_cast_808_wire_constant <= "00000000000000000000000000000010";
    type_cast_814_wire_constant <= "00000000000000000000000000000001";
    type_cast_820_wire_constant <= "11111111111111111111111111111111";
    type_cast_830_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_837_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_846_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_860_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_865_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_93_wire_constant <= "00000000000000000000000000001000";
    type_cast_947_wire_constant <= "00000000";
    type_cast_951_wire_constant <= "00000000";
    type_cast_955_wire_constant <= "00000000";
    type_cast_959_wire_constant <= "00000000";
    phi_stmt_1340: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1344_wire_constant & type_cast_1346_wire;
      req <= phi_stmt_1340_req_0 & phi_stmt_1340_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1340",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1340_ack_0,
          idata => idata,
          odata => indvar_1340,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1340
    phi_stmt_403: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_407_wire_constant & type_cast_409_wire;
      req <= phi_stmt_403_req_0 & phi_stmt_403_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_403",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_403_ack_0,
          idata => idata,
          odata => indvar795_403,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_403
    phi_stmt_610: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_614_wire_constant & type_cast_616_wire;
      req <= phi_stmt_610_req_0 & phi_stmt_610_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_610",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_610_ack_0,
          idata => idata,
          odata => indvar783_610,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_610
    phi_stmt_842: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_846_wire_constant & type_cast_848_wire;
      req <= phi_stmt_842_req_0 & phi_stmt_842_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_842",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_842_ack_0,
          idata => idata,
          odata => indvar772_842,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_842
    -- flow-through select operator MUX_1336_inst
    tmp771_1337 <= xx_xop_1330 when (tmp768_1314(0) /=  '0') else type_cast_1335_wire_constant;
    -- flow-through select operator MUX_399_inst
    tmp804_400 <= xx_xop808_393 when (tmp800_377(0) /=  '0') else type_cast_398_wire_constant;
    -- flow-through select operator MUX_606_inst
    tmp793_607 <= xx_xop807_600 when (tmp789_584(0) /=  '0') else type_cast_605_wire_constant;
    -- flow-through select operator MUX_838_inst
    tmp781_839 <= xx_xop806_832 when (tmp777_816(0) /=  '0') else type_cast_837_wire_constant;
    addr_of_1353_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1353_final_reg_req_0;
      addr_of_1353_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1353_final_reg_req_1;
      addr_of_1353_final_reg_ack_1<= rack(0);
      addr_of_1353_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1353_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1352_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx635_1354,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_416_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_416_final_reg_req_0;
      addr_of_416_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_416_final_reg_req_1;
      addr_of_416_final_reg_ack_1<= rack(0);
      addr_of_416_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_416_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_415_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_623_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_623_final_reg_req_0;
      addr_of_623_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_623_final_reg_req_1;
      addr_of_623_final_reg_ack_1<= rack(0);
      addr_of_623_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_623_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_622_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_624,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_855_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_855_final_reg_req_0;
      addr_of_855_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_855_final_reg_req_1;
      addr_of_855_final_reg_ack_1<= rack(0);
      addr_of_855_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_855_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_854_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_856,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_101_inst_req_0;
      type_cast_101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_101_inst_req_1;
      type_cast_101_inst_ack_1<= rack(0);
      type_cast_101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1035_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1035_inst_req_0;
      type_cast_1035_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1035_inst_req_1;
      type_cast_1035_inst_ack_1<= rack(0);
      type_cast_1035_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1035_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv415_1036,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1048_inst_req_0;
      type_cast_1048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1048_inst_req_1;
      type_cast_1048_inst_ack_1<= rack(0);
      type_cast_1048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr417_1045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv418_1049,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1143_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1143_inst_req_0;
      type_cast_1143_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1143_inst_req_1;
      type_cast_1143_inst_ack_1<= rack(0);
      type_cast_1143_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1143_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr500_1140,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv501_1144,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr583_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv584_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1285_inst_req_0;
      type_cast_1285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1285_inst_req_1;
      type_cast_1285_inst_ack_1<= rack(0);
      type_cast_1285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1284_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv619_1286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1323_inst_req_0;
      type_cast_1323_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1323_inst_req_1;
      type_cast_1323_inst_ack_1<= rack(0);
      type_cast_1323_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1323_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp767x_xop_1320,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_292_1324,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1346_inst_req_0;
      type_cast_1346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1346_inst_req_1;
      type_cast_1346_inst_ack_1<= rack(0);
      type_cast_1346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1346_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1361_inst_req_0;
      type_cast_1361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1361_inst_req_1;
      type_cast_1361_inst_ack_1<= rack(0);
      type_cast_1361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp636_1358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv639_1362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1371_inst_req_0;
      type_cast_1371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1371_inst_req_1;
      type_cast_1371_inst_ack_1<= rack(0);
      type_cast_1371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1371_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr642_1368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv645_1372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1381_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1381_inst_req_0;
      type_cast_1381_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1381_inst_req_1;
      type_cast_1381_inst_ack_1<= rack(0);
      type_cast_1381_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1381_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr648_1378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv651_1382,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_138_inst_req_0;
      type_cast_138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_138_inst_req_1;
      type_cast_138_inst_ack_1<= rack(0);
      type_cast_138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1391_inst_req_0;
      type_cast_1391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1391_inst_req_1;
      type_cast_1391_inst_ack_1<= rack(0);
      type_cast_1391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr654_1388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv657_1392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1401_inst_req_0;
      type_cast_1401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1401_inst_req_1;
      type_cast_1401_inst_ack_1<= rack(0);
      type_cast_1401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr660_1398,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv663_1402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1411_inst_req_0;
      type_cast_1411_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1411_inst_req_1;
      type_cast_1411_inst_ack_1<= rack(0);
      type_cast_1411_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1411_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr666_1408,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv669_1412,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1421_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1421_inst_req_0;
      type_cast_1421_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1421_inst_req_1;
      type_cast_1421_inst_ack_1<= rack(0);
      type_cast_1421_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1421_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr672_1418,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv675_1422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1431_inst_req_0;
      type_cast_1431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1431_inst_req_1;
      type_cast_1431_inst_ack_1<= rack(0);
      type_cast_1431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr678_1428,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv681_1432,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_151_inst_req_0;
      type_cast_151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_151_inst_req_1;
      type_cast_151_inst_ack_1<= rack(0);
      type_cast_151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_163_inst_req_0;
      type_cast_163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_163_inst_req_1;
      type_cast_163_inst_ack_1<= rack(0);
      type_cast_163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_176_inst_req_0;
      type_cast_176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_176_inst_req_1;
      type_cast_176_inst_ack_1<= rack(0);
      type_cast_176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_188_inst_req_0;
      type_cast_188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_188_inst_req_1;
      type_cast_188_inst_ack_1<= rack(0);
      type_cast_188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_201_inst_req_0;
      type_cast_201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_201_inst_req_1;
      type_cast_201_inst_ack_1<= rack(0);
      type_cast_201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_273_inst_req_0;
      type_cast_273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_273_inst_req_1;
      type_cast_273_inst_ack_1<= rack(0);
      type_cast_273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_270,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_286_inst_req_0;
      type_cast_286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_286_inst_req_1;
      type_cast_286_inst_ack_1<= rack(0);
      type_cast_286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_283,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_298_inst_req_0;
      type_cast_298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_298_inst_req_1;
      type_cast_298_inst_ack_1<= rack(0);
      type_cast_298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_295,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_311_inst_req_0;
      type_cast_311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_311_inst_req_1;
      type_cast_311_inst_ack_1<= rack(0);
      type_cast_311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_312,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_323_inst_req_0;
      type_cast_323_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_323_inst_req_1;
      type_cast_323_inst_ack_1<= rack(0);
      type_cast_323_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_323_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_320,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_324,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_336_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_336_inst_req_0;
      type_cast_336_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_336_inst_req_1;
      type_cast_336_inst_ack_1<= rack(0);
      type_cast_336_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_336_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_333,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_337,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_386_inst_req_0;
      type_cast_386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_386_inst_req_1;
      type_cast_386_inst_ack_1<= rack(0);
      type_cast_386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp799x_xop_383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_387,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_409_inst_req_0;
      type_cast_409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_409_inst_req_1;
      type_cast_409_inst_ack_1<= rack(0);
      type_cast_409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext796_560,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_409_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_423_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_423_inst_req_0;
      type_cast_423_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_423_inst_req_1;
      type_cast_423_inst_ack_1<= rack(0);
      type_cast_423_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_423_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_424,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_436_inst_req_0;
      type_cast_436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_436_inst_req_1;
      type_cast_436_inst_ack_1<= rack(0);
      type_cast_436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_433,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_437,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_454_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_454_inst_req_0;
      type_cast_454_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_454_inst_req_1;
      type_cast_454_inst_ack_1<= rack(0);
      type_cast_454_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_454_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_451,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_455,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_472_inst_req_0;
      type_cast_472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_472_inst_req_1;
      type_cast_472_inst_ack_1<= rack(0);
      type_cast_472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_469,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_490_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_490_inst_req_0;
      type_cast_490_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_490_inst_req_1;
      type_cast_490_inst_ack_1<= rack(0);
      type_cast_490_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_490_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_491,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_508_inst_req_0;
      type_cast_508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_508_inst_req_1;
      type_cast_508_inst_ack_1<= rack(0);
      type_cast_508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_505,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_51_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_51_inst_req_0;
      type_cast_51_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_51_inst_req_1;
      type_cast_51_inst_ack_1<= rack(0);
      type_cast_51_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_51_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_48,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_52,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_526_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_526_inst_req_0;
      type_cast_526_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_526_inst_req_1;
      type_cast_526_inst_ack_1<= rack(0);
      type_cast_526_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_526_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_523,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_527,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_544_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_544_inst_req_0;
      type_cast_544_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_544_inst_req_1;
      type_cast_544_inst_ack_1<= rack(0);
      type_cast_544_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_544_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_541,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_545,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_593_inst_req_0;
      type_cast_593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_593_inst_req_1;
      type_cast_593_inst_ack_1<= rack(0);
      type_cast_593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_593_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp788x_xop_590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_594,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_616_inst_req_0;
      type_cast_616_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_616_inst_req_1;
      type_cast_616_inst_ack_1<= rack(0);
      type_cast_616_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_616_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext784_767,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_616_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_630_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_630_inst_req_0;
      type_cast_630_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_630_inst_req_1;
      type_cast_630_inst_ack_1<= rack(0);
      type_cast_630_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_630_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_643_inst_req_0;
      type_cast_643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_643_inst_req_1;
      type_cast_643_inst_ack_1<= rack(0);
      type_cast_643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_643_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_640,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_661_inst_req_0;
      type_cast_661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_661_inst_req_1;
      type_cast_661_inst_ack_1<= rack(0);
      type_cast_661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_662,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_679_inst_req_0;
      type_cast_679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_679_inst_req_1;
      type_cast_679_inst_ack_1<= rack(0);
      type_cast_679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_680,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_697_inst_req_0;
      type_cast_697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_697_inst_req_1;
      type_cast_697_inst_ack_1<= rack(0);
      type_cast_697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_694,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_715_inst_req_0;
      type_cast_715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_715_inst_req_1;
      type_cast_715_inst_ack_1<= rack(0);
      type_cast_715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_712,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_733_inst_req_0;
      type_cast_733_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_733_inst_req_1;
      type_cast_733_inst_ack_1<= rack(0);
      type_cast_733_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_733_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_730,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_734,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_751_inst_req_0;
      type_cast_751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_751_inst_req_1;
      type_cast_751_inst_ack_1<= rack(0);
      type_cast_751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_825_inst_req_0;
      type_cast_825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_825_inst_req_1;
      type_cast_825_inst_ack_1<= rack(0);
      type_cast_825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp776x_xop_822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_848_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_848_inst_req_0;
      type_cast_848_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_848_inst_req_1;
      type_cast_848_inst_ack_1<= rack(0);
      type_cast_848_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_848_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext773_867,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_848_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_889_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_889_inst_req_0;
      type_cast_889_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_889_inst_req_1;
      type_cast_889_inst_ack_1<= rack(0);
      type_cast_889_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_889_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_888_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_890,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1352_index_1_rename
    process(R_indvar_1351_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1351_resized;
      ov(13 downto 0) := iv;
      R_indvar_1351_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1352_index_1_resize
    process(indvar_1340) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1340;
      ov := iv(13 downto 0);
      R_indvar_1351_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1352_root_address_inst
    process(array_obj_ref_1352_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1352_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1352_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_415_index_1_rename
    process(R_indvar795_414_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar795_414_resized;
      ov(13 downto 0) := iv;
      R_indvar795_414_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_415_index_1_resize
    process(indvar795_403) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar795_403;
      ov := iv(13 downto 0);
      R_indvar795_414_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_415_root_address_inst
    process(array_obj_ref_415_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_415_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_415_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_622_index_1_rename
    process(R_indvar783_621_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar783_621_resized;
      ov(10 downto 0) := iv;
      R_indvar783_621_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_622_index_1_resize
    process(indvar783_610) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar783_610;
      ov := iv(10 downto 0);
      R_indvar783_621_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_622_root_address_inst
    process(array_obj_ref_622_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_622_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_622_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_854_index_1_rename
    process(R_indvar772_853_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar772_853_resized;
      ov(13 downto 0) := iv;
      R_indvar772_853_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_854_index_1_resize
    process(indvar772_842) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar772_842;
      ov := iv(13 downto 0);
      R_indvar772_853_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_854_root_address_inst
    process(array_obj_ref_854_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_854_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_854_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1357_addr_0
    process(ptr_deref_1357_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1357_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1357_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1357_base_resize
    process(arrayidx635_1354) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx635_1354;
      ov := iv(13 downto 0);
      ptr_deref_1357_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1357_gather_scatter
    process(ptr_deref_1357_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1357_data_0;
      ov(63 downto 0) := iv;
      tmp636_1358 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1357_root_address_inst
    process(ptr_deref_1357_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1357_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1357_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_552_addr_0
    process(ptr_deref_552_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_552_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_552_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_552_base_resize
    process(arrayidx_417) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_417;
      ov := iv(13 downto 0);
      ptr_deref_552_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_552_gather_scatter
    process(add186_550) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_550;
      ov(63 downto 0) := iv;
      ptr_deref_552_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_552_root_address_inst
    process(ptr_deref_552_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_552_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_552_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_759_addr_0
    process(ptr_deref_759_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_759_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_759_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_759_base_resize
    process(arrayidx246_624) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_624;
      ov := iv(10 downto 0);
      ptr_deref_759_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_759_gather_scatter
    process(add242_757) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_757;
      ov(63 downto 0) := iv;
      ptr_deref_759_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_759_root_address_inst
    process(ptr_deref_759_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_759_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_759_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_858_addr_0
    process(ptr_deref_858_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_858_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_858_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_858_base_resize
    process(arrayidx269_856) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_856;
      ov := iv(13 downto 0);
      ptr_deref_858_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_858_gather_scatter
    process(type_cast_860_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_860_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_858_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_858_root_address_inst
    process(ptr_deref_858_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_858_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_858_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1296_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264755_797;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1296_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1296_branch_req_0,
          ack0 => if_stmt_1296_branch_ack_0,
          ack1 => if_stmt_1296_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1468_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1467;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1468_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1468_branch_req_0,
          ack0 => if_stmt_1468_branch_ack_0,
          ack1 => if_stmt_1468_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_350_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp763_349;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_350_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_350_branch_req_0,
          ack0 => if_stmt_350_branch_ack_0,
          ack1 => if_stmt_350_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_365_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194759_364;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_365_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_365_branch_req_0,
          ack0 => if_stmt_365_branch_ack_0,
          ack1 => if_stmt_365_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_566_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_565;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_566_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_566_branch_req_0,
          ack0 => if_stmt_566_branch_ack_0,
          ack1 => if_stmt_566_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_773_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_772;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_773_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_773_branch_req_0,
          ack0 => if_stmt_773_branch_ack_0,
          ack1 => if_stmt_773_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_798_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264755_797;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_798_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_798_branch_req_0,
          ack0 => if_stmt_798_branch_ack_0,
          ack1 => if_stmt_798_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_873_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_872;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_873_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_873_branch_req_0,
          ack0 => if_stmt_873_branch_ack_0,
          ack1 => if_stmt_873_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1319_inst
    process(tmp767_1308) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp767_1308, type_cast_1318_wire_constant, tmp_var);
      tmp767x_xop_1320 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_239_inst
    process(add74_235, shr_223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_235, shr_223, tmp_var);
      add79_240 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_382_inst
    process(shr_223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_223, type_cast_381_wire_constant, tmp_var);
      tmp799x_xop_383 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_589_inst
    process(tmp788_578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp788_578, type_cast_588_wire_constant, tmp_var);
      tmp788x_xop_590 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_821_inst
    process(tmp776_810) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp776_810, type_cast_820_wire_constant, tmp_var);
      tmp776x_xop_822 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1329_inst
    process(iNsTr_292_1324) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_292_1324, type_cast_1328_wire_constant, tmp_var);
      xx_xop_1330 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1461_inst
    process(indvar_1340) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1340, type_cast_1460_wire_constant, tmp_var);
      indvarx_xnext_1462 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_392_inst
    process(iNsTr_26_387) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_387, type_cast_391_wire_constant, tmp_var);
      xx_xop808_393 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_559_inst
    process(indvar795_403) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar795_403, type_cast_558_wire_constant, tmp_var);
      indvarx_xnext796_560 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_599_inst
    process(iNsTr_39_594) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_594, type_cast_598_wire_constant, tmp_var);
      xx_xop807_600 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_766_inst
    process(indvar783_610) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar783_610, type_cast_765_wire_constant, tmp_var);
      indvarx_xnext784_767 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_831_inst
    process(iNsTr_53_826) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_826, type_cast_830_wire_constant, tmp_var);
      xx_xop806_832 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_866_inst
    process(indvar772_842) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar772_842, type_cast_865_wire_constant, tmp_var);
      indvarx_xnext773_867 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_234_inst
    process(iNsTr_14_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_229, type_cast_233_wire_constant, tmp_var);
      add74_235 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1466_inst
    process(indvarx_xnext_1462, tmp771_1337) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1462, tmp771_1337, tmp_var);
      exitcond1_1467 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_564_inst
    process(indvarx_xnext796_560, tmp804_400) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext796_560, tmp804_400, tmp_var);
      exitcond3_565 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_771_inst
    process(indvarx_xnext784_767, tmp793_607) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext784_767, tmp793_607, tmp_var);
      exitcond2_772 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_871_inst
    process(indvarx_xnext773_867, tmp781_839) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext773_867, tmp781_839, tmp_var);
      exitcond_872 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1044_inst
    process(mul66_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_217, type_cast_1043_wire_constant, tmp_var);
      shr417_1045 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1139_inst
    process(mul66_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_217, type_cast_1138_wire_constant, tmp_var);
      shr500_1140 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1234_inst
    process(add79_240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_240, type_cast_1233_wire_constant, tmp_var);
      shr583_1235 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1307_inst
    process(mul259_791) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_791, type_cast_1306_wire_constant, tmp_var);
      tmp767_1308 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_222_inst
    process(mul66_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_217, type_cast_221_wire_constant, tmp_var);
      shr_223 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_228_inst
    process(mul66_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_217, type_cast_227_wire_constant, tmp_var);
      iNsTr_14_229 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_577_inst
    process(mul91_255) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_255, type_cast_576_wire_constant, tmp_var);
      tmp788_578 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_809_inst
    process(mul259_791) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_791, type_cast_808_wire_constant, tmp_var);
      tmp776_810 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1367_inst
    process(tmp636_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp636_1358, type_cast_1366_wire_constant, tmp_var);
      shr642_1368 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1377_inst
    process(tmp636_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp636_1358, type_cast_1376_wire_constant, tmp_var);
      shr648_1378 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1387_inst
    process(tmp636_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp636_1358, type_cast_1386_wire_constant, tmp_var);
      shr654_1388 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1397_inst
    process(tmp636_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp636_1358, type_cast_1396_wire_constant, tmp_var);
      shr660_1398 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1407_inst
    process(tmp636_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp636_1358, type_cast_1406_wire_constant, tmp_var);
      shr666_1408 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1417_inst
    process(tmp636_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp636_1358, type_cast_1416_wire_constant, tmp_var);
      shr672_1418 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1427_inst
    process(tmp636_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp636_1358, type_cast_1426_wire_constant, tmp_var);
      shr678_1428 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_211_inst
    process(add12_82, add_57) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add12_82, add_57, tmp_var);
      mul_212 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_216_inst
    process(mul_212, add21_107) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_212, add21_107, tmp_var);
      mul66_217 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_244_inst
    process(add39_157, add30_132) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add39_157, add30_132, tmp_var);
      mul85_245 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_249_inst
    process(mul85_245, add48_182) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_245, add48_182, tmp_var);
      mul88_250 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_254_inst
    process(mul88_250, add57_207) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_250, add57_207, tmp_var);
      mul91_255 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_785_inst
    process(add126_317, add117_292) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add126_317, add117_292, tmp_var);
      mul256_786 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_790_inst
    process(mul256_786, add135_342) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_786, add135_342, tmp_var);
      mul259_791 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_106_inst
    process(shl18_95, conv20_102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_95, conv20_102, tmp_var);
      add21_107 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_131_inst
    process(shl27_120, conv29_127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_120, conv29_127, tmp_var);
      add30_132 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_156_inst
    process(shl36_145, conv38_152) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_145, conv38_152, tmp_var);
      add39_157 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_181_inst
    process(shl45_170, conv47_177) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_170, conv47_177, tmp_var);
      add48_182 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_206_inst
    process(shl54_195, conv56_202) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_195, conv56_202, tmp_var);
      add57_207 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_291_inst
    process(shl114_280, conv116_287) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_280, conv116_287, tmp_var);
      add117_292 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_316_inst
    process(shl123_305, conv125_312) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_305, conv125_312, tmp_var);
      add126_317 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_341_inst
    process(shl132_330, conv134_337) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_330, conv134_337, tmp_var);
      add135_342 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_56_inst
    process(shl_45, conv3_52) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_45, conv3_52, tmp_var);
      add_57 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_81_inst
    process(shl9_70, conv11_77) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_70, conv11_77, tmp_var);
      add12_82 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_441_inst
    process(shl146_430, conv149_437) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_430, conv149_437, tmp_var);
      add150_442 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_459_inst
    process(shl152_448, conv155_455) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_448, conv155_455, tmp_var);
      add156_460 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_477_inst
    process(shl158_466, conv161_473) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_466, conv161_473, tmp_var);
      add162_478 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_495_inst
    process(shl164_484, conv167_491) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_484, conv167_491, tmp_var);
      add168_496 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_513_inst
    process(shl170_502, conv173_509) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_502, conv173_509, tmp_var);
      add174_514 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_531_inst
    process(shl176_520, conv179_527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_520, conv179_527, tmp_var);
      add180_532 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_549_inst
    process(shl182_538, conv185_545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_538, conv185_545, tmp_var);
      add186_550 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_648_inst
    process(shl202_637, conv205_644) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_637, conv205_644, tmp_var);
      add206_649 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_666_inst
    process(shl208_655, conv211_662) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_655, conv211_662, tmp_var);
      add212_667 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_684_inst
    process(shl214_673, conv217_680) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_673, conv217_680, tmp_var);
      add218_685 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_702_inst
    process(shl220_691, conv223_698) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_691, conv223_698, tmp_var);
      add224_703 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_720_inst
    process(shl226_709, conv229_716) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_709, conv229_716, tmp_var);
      add230_721 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_738_inst
    process(shl232_727, conv235_734) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_727, conv235_734, tmp_var);
      add236_739 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_756_inst
    process(shl238_745, conv241_752) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_745, conv241_752, tmp_var);
      add242_757 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_119_inst
    process(conv26_114) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_114, type_cast_118_wire_constant, tmp_var);
      shl27_120 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_144_inst
    process(conv35_139) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_139, type_cast_143_wire_constant, tmp_var);
      shl36_145 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_169_inst
    process(conv44_164) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_164, type_cast_168_wire_constant, tmp_var);
      shl45_170 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_194_inst
    process(conv53_189) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_189, type_cast_193_wire_constant, tmp_var);
      shl54_195 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_279_inst
    process(conv113_274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_274, type_cast_278_wire_constant, tmp_var);
      shl114_280 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_304_inst
    process(conv122_299) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_299, type_cast_303_wire_constant, tmp_var);
      shl123_305 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_329_inst
    process(conv131_324) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_324, type_cast_328_wire_constant, tmp_var);
      shl132_330 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_44_inst
    process(conv1_39) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_39, type_cast_43_wire_constant, tmp_var);
      shl_45 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_69_inst
    process(conv8_64) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_64, type_cast_68_wire_constant, tmp_var);
      shl9_70 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_94_inst
    process(conv17_89) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_89, type_cast_93_wire_constant, tmp_var);
      shl18_95 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_429_inst
    process(conv144_424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_424, type_cast_428_wire_constant, tmp_var);
      shl146_430 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_447_inst
    process(add150_442) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_442, type_cast_446_wire_constant, tmp_var);
      shl152_448 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_465_inst
    process(add156_460) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_460, type_cast_464_wire_constant, tmp_var);
      shl158_466 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_483_inst
    process(add162_478) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_478, type_cast_482_wire_constant, tmp_var);
      shl164_484 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_501_inst
    process(add168_496) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_496, type_cast_500_wire_constant, tmp_var);
      shl170_502 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_519_inst
    process(add174_514) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_514, type_cast_518_wire_constant, tmp_var);
      shl176_520 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_537_inst
    process(add180_532) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_532, type_cast_536_wire_constant, tmp_var);
      shl182_538 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_636_inst
    process(conv200_631) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_631, type_cast_635_wire_constant, tmp_var);
      shl202_637 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_654_inst
    process(add206_649) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_649, type_cast_653_wire_constant, tmp_var);
      shl208_655 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_672_inst
    process(add212_667) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_667, type_cast_671_wire_constant, tmp_var);
      shl214_673 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_690_inst
    process(add218_685) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_685, type_cast_689_wire_constant, tmp_var);
      shl220_691 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_708_inst
    process(add224_703) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_703, type_cast_707_wire_constant, tmp_var);
      shl226_709 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_726_inst
    process(add230_721) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_721, type_cast_725_wire_constant, tmp_var);
      shl232_727 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_744_inst
    process(add236_739) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_739, type_cast_743_wire_constant, tmp_var);
      shl238_745 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1290_inst
    process(conv619_1286, conv276_890) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv619_1286, conv276_890, tmp_var);
      sub_1291 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1313_inst
    process(tmp767_1308) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp767_1308, type_cast_1312_wire_constant, tmp_var);
      tmp768_1314 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_347_inst
    process(mul66_217) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_217, type_cast_346_wire_constant, tmp_var);
      cmp763_349 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_363_inst
    process(mul91_255) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_255, type_cast_362_wire_constant, tmp_var);
      cmp194759_364 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_376_inst
    process(shr_223) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_223, type_cast_375_wire_constant, tmp_var);
      tmp800_377 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_583_inst
    process(tmp788_578) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp788_578, type_cast_582_wire_constant, tmp_var);
      tmp789_584 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_796_inst
    process(mul259_791) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_791, type_cast_795_wire_constant, tmp_var);
      cmp264755_797 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_815_inst
    process(tmp776_810) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp776_810, type_cast_814_wire_constant, tmp_var);
      tmp777_816 <= tmp_var; --
    end process;
    -- shared split operator group (96) : array_obj_ref_1352_index_offset 
    ApIntAdd_group_96: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1351_scaled;
      array_obj_ref_1352_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1352_index_offset_req_0;
      array_obj_ref_1352_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1352_index_offset_req_1;
      array_obj_ref_1352_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_96_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_96_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_96",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 96
    -- shared split operator group (97) : array_obj_ref_415_index_offset 
    ApIntAdd_group_97: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar795_414_scaled;
      array_obj_ref_415_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_415_index_offset_req_0;
      array_obj_ref_415_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_415_index_offset_req_1;
      array_obj_ref_415_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_97_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_97_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_97",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 97
    -- shared split operator group (98) : array_obj_ref_622_index_offset 
    ApIntAdd_group_98: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar783_621_scaled;
      array_obj_ref_622_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_622_index_offset_req_0;
      array_obj_ref_622_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_622_index_offset_req_1;
      array_obj_ref_622_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_98_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_98_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_98",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 98
    -- shared split operator group (99) : array_obj_ref_854_index_offset 
    ApIntAdd_group_99: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar772_853_scaled;
      array_obj_ref_854_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_854_index_offset_req_0;
      array_obj_ref_854_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_854_index_offset_req_1;
      array_obj_ref_854_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_99_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_99_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_99",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 99
    -- unary operator type_cast_1284_inst
    process(call618_1281) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call618_1281, tmp_var);
      type_cast_1284_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_888_inst
    process(call275_884) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_884, tmp_var);
      type_cast_888_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1357_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1357_load_0_req_0;
      ptr_deref_1357_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1357_load_0_req_1;
      ptr_deref_1357_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1357_word_address_0;
      ptr_deref_1357_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_552_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_552_store_0_req_0;
      ptr_deref_552_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_552_store_0_req_1;
      ptr_deref_552_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_552_word_address_0;
      data_in <= ptr_deref_552_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_759_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_759_store_0_req_0;
      ptr_deref_759_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_759_store_0_req_1;
      ptr_deref_759_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_759_word_address_0;
      data_in <= ptr_deref_759_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_858_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_858_store_0_req_0;
      ptr_deref_858_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_858_store_0_req_1;
      ptr_deref_858_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_858_word_address_0;
      data_in <= ptr_deref_858_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1268_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1268_inst_req_0;
      RPIPE_Block0_done_1268_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1268_inst_req_1;
      RPIPE_Block0_done_1268_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call610_1269 <= data_out(7 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1271_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1271_inst_req_0;
      RPIPE_Block1_done_1271_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1271_inst_req_1;
      RPIPE_Block1_done_1271_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call612_1272 <= data_out(7 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1274_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1274_inst_req_0;
      RPIPE_Block2_done_1274_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1274_inst_req_1;
      RPIPE_Block2_done_1274_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call614_1275 <= data_out(7 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1277_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1277_inst_req_0;
      RPIPE_Block3_done_1277_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1277_inst_req_1;
      RPIPE_Block3_done_1277_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call616_1278 <= data_out(7 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_47_inst RPIPE_ConvTranspose_input_pipe_59_inst RPIPE_ConvTranspose_input_pipe_72_inst RPIPE_ConvTranspose_input_pipe_84_inst RPIPE_ConvTranspose_input_pipe_97_inst RPIPE_ConvTranspose_input_pipe_109_inst RPIPE_ConvTranspose_input_pipe_122_inst RPIPE_ConvTranspose_input_pipe_134_inst RPIPE_ConvTranspose_input_pipe_147_inst RPIPE_ConvTranspose_input_pipe_159_inst RPIPE_ConvTranspose_input_pipe_172_inst RPIPE_ConvTranspose_input_pipe_184_inst RPIPE_ConvTranspose_input_pipe_197_inst RPIPE_ConvTranspose_input_pipe_257_inst RPIPE_ConvTranspose_input_pipe_260_inst RPIPE_ConvTranspose_input_pipe_263_inst RPIPE_ConvTranspose_input_pipe_266_inst RPIPE_ConvTranspose_input_pipe_269_inst RPIPE_ConvTranspose_input_pipe_282_inst RPIPE_ConvTranspose_input_pipe_294_inst RPIPE_ConvTranspose_input_pipe_307_inst RPIPE_ConvTranspose_input_pipe_319_inst RPIPE_ConvTranspose_input_pipe_332_inst RPIPE_ConvTranspose_input_pipe_419_inst RPIPE_ConvTranspose_input_pipe_432_inst RPIPE_ConvTranspose_input_pipe_450_inst RPIPE_ConvTranspose_input_pipe_468_inst RPIPE_ConvTranspose_input_pipe_486_inst RPIPE_ConvTranspose_input_pipe_504_inst RPIPE_ConvTranspose_input_pipe_522_inst RPIPE_ConvTranspose_input_pipe_540_inst RPIPE_ConvTranspose_input_pipe_626_inst RPIPE_ConvTranspose_input_pipe_639_inst RPIPE_ConvTranspose_input_pipe_657_inst RPIPE_ConvTranspose_input_pipe_675_inst RPIPE_ConvTranspose_input_pipe_693_inst RPIPE_ConvTranspose_input_pipe_711_inst RPIPE_ConvTranspose_input_pipe_729_inst RPIPE_ConvTranspose_input_pipe_747_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_257_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_260_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_263_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_266_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_269_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_282_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_294_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_307_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_319_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_332_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_419_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_432_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_450_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_468_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_486_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_504_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_522_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_540_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_626_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_639_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_657_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_675_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_693_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_711_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_729_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_747_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_257_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_260_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_263_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_266_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_269_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_282_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_294_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_307_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_319_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_332_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_419_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_432_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_450_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_468_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_486_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_504_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_522_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_540_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_626_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_639_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_657_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_675_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_693_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_711_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_729_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_747_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_257_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_260_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_263_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_266_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_269_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_282_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_294_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_307_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_319_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_332_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_419_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_432_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_450_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_468_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_486_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_504_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_522_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_540_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_626_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_639_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_657_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_675_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_693_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_711_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_729_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_747_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_257_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_260_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_263_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_266_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_269_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_282_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_294_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_307_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_319_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_332_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_419_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_432_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_450_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_468_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_486_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_504_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_522_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_540_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_626_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_639_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_657_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_675_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_693_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_711_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_729_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_747_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call_35 <= data_out(319 downto 312);
      call2_48 <= data_out(311 downto 304);
      call5_60 <= data_out(303 downto 296);
      call10_73 <= data_out(295 downto 288);
      call14_85 <= data_out(287 downto 280);
      call19_98 <= data_out(279 downto 272);
      call23_110 <= data_out(271 downto 264);
      call28_123 <= data_out(263 downto 256);
      call32_135 <= data_out(255 downto 248);
      call37_148 <= data_out(247 downto 240);
      call41_160 <= data_out(239 downto 232);
      call46_173 <= data_out(231 downto 224);
      call50_185 <= data_out(223 downto 216);
      call55_198 <= data_out(215 downto 208);
      call92_258 <= data_out(207 downto 200);
      call97_261 <= data_out(199 downto 192);
      call101_264 <= data_out(191 downto 184);
      call106_267 <= data_out(183 downto 176);
      call110_270 <= data_out(175 downto 168);
      call115_283 <= data_out(167 downto 160);
      call119_295 <= data_out(159 downto 152);
      call124_308 <= data_out(151 downto 144);
      call128_320 <= data_out(143 downto 136);
      call133_333 <= data_out(135 downto 128);
      call143_420 <= data_out(127 downto 120);
      call147_433 <= data_out(119 downto 112);
      call153_451 <= data_out(111 downto 104);
      call159_469 <= data_out(103 downto 96);
      call165_487 <= data_out(95 downto 88);
      call171_505 <= data_out(87 downto 80);
      call177_523 <= data_out(79 downto 72);
      call183_541 <= data_out(71 downto 64);
      call199_627 <= data_out(63 downto 56);
      call203_640 <= data_out(55 downto 48);
      call209_658 <= data_out(47 downto 40);
      call215_676 <= data_out(39 downto 32);
      call221_694 <= data_out(31 downto 24);
      call227_712 <= data_out(23 downto 16);
      call233_730 <= data_out(15 downto 8);
      call239_748 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_894_inst WPIPE_Block0_start_936_inst WPIPE_Block0_start_897_inst WPIPE_Block0_start_921_inst WPIPE_Block0_start_903_inst WPIPE_Block0_start_939_inst WPIPE_Block0_start_927_inst WPIPE_Block0_start_942_inst WPIPE_Block0_start_945_inst WPIPE_Block0_start_949_inst WPIPE_Block0_start_906_inst WPIPE_Block0_start_953_inst WPIPE_Block0_start_930_inst WPIPE_Block0_start_957_inst WPIPE_Block0_start_909_inst WPIPE_Block0_start_912_inst WPIPE_Block0_start_933_inst WPIPE_Block0_start_961_inst WPIPE_Block0_start_964_inst WPIPE_Block0_start_915_inst WPIPE_Block0_start_967_inst WPIPE_Block0_start_970_inst WPIPE_Block0_start_918_inst WPIPE_Block0_start_973_inst WPIPE_Block0_start_976_inst WPIPE_Block0_start_924_inst WPIPE_Block0_start_900_inst WPIPE_Block0_start_891_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 27 downto 0);
      signal update_req, update_ack : BooleanArray( 27 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 27 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant inBUFs : IntegerArray(27 downto 0) := (27 => 0, 26 => 0, 25 => 0, 24 => 0, 23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      sample_req_unguarded(27) <= WPIPE_Block0_start_894_inst_req_0;
      sample_req_unguarded(26) <= WPIPE_Block0_start_936_inst_req_0;
      sample_req_unguarded(25) <= WPIPE_Block0_start_897_inst_req_0;
      sample_req_unguarded(24) <= WPIPE_Block0_start_921_inst_req_0;
      sample_req_unguarded(23) <= WPIPE_Block0_start_903_inst_req_0;
      sample_req_unguarded(22) <= WPIPE_Block0_start_939_inst_req_0;
      sample_req_unguarded(21) <= WPIPE_Block0_start_927_inst_req_0;
      sample_req_unguarded(20) <= WPIPE_Block0_start_942_inst_req_0;
      sample_req_unguarded(19) <= WPIPE_Block0_start_945_inst_req_0;
      sample_req_unguarded(18) <= WPIPE_Block0_start_949_inst_req_0;
      sample_req_unguarded(17) <= WPIPE_Block0_start_906_inst_req_0;
      sample_req_unguarded(16) <= WPIPE_Block0_start_953_inst_req_0;
      sample_req_unguarded(15) <= WPIPE_Block0_start_930_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Block0_start_957_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Block0_start_909_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_912_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_933_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_961_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_964_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_915_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_967_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_970_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_918_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_973_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_976_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_924_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_900_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_891_inst_req_0;
      WPIPE_Block0_start_894_inst_ack_0 <= sample_ack_unguarded(27);
      WPIPE_Block0_start_936_inst_ack_0 <= sample_ack_unguarded(26);
      WPIPE_Block0_start_897_inst_ack_0 <= sample_ack_unguarded(25);
      WPIPE_Block0_start_921_inst_ack_0 <= sample_ack_unguarded(24);
      WPIPE_Block0_start_903_inst_ack_0 <= sample_ack_unguarded(23);
      WPIPE_Block0_start_939_inst_ack_0 <= sample_ack_unguarded(22);
      WPIPE_Block0_start_927_inst_ack_0 <= sample_ack_unguarded(21);
      WPIPE_Block0_start_942_inst_ack_0 <= sample_ack_unguarded(20);
      WPIPE_Block0_start_945_inst_ack_0 <= sample_ack_unguarded(19);
      WPIPE_Block0_start_949_inst_ack_0 <= sample_ack_unguarded(18);
      WPIPE_Block0_start_906_inst_ack_0 <= sample_ack_unguarded(17);
      WPIPE_Block0_start_953_inst_ack_0 <= sample_ack_unguarded(16);
      WPIPE_Block0_start_930_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Block0_start_957_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Block0_start_909_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_912_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_933_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_961_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_964_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_915_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_967_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_970_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_918_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_973_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_976_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_924_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_900_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_891_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(27) <= WPIPE_Block0_start_894_inst_req_1;
      update_req_unguarded(26) <= WPIPE_Block0_start_936_inst_req_1;
      update_req_unguarded(25) <= WPIPE_Block0_start_897_inst_req_1;
      update_req_unguarded(24) <= WPIPE_Block0_start_921_inst_req_1;
      update_req_unguarded(23) <= WPIPE_Block0_start_903_inst_req_1;
      update_req_unguarded(22) <= WPIPE_Block0_start_939_inst_req_1;
      update_req_unguarded(21) <= WPIPE_Block0_start_927_inst_req_1;
      update_req_unguarded(20) <= WPIPE_Block0_start_942_inst_req_1;
      update_req_unguarded(19) <= WPIPE_Block0_start_945_inst_req_1;
      update_req_unguarded(18) <= WPIPE_Block0_start_949_inst_req_1;
      update_req_unguarded(17) <= WPIPE_Block0_start_906_inst_req_1;
      update_req_unguarded(16) <= WPIPE_Block0_start_953_inst_req_1;
      update_req_unguarded(15) <= WPIPE_Block0_start_930_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Block0_start_957_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Block0_start_909_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_912_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_933_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_961_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_964_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_915_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_967_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_970_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_918_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_973_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_976_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_924_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_900_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_891_inst_req_1;
      WPIPE_Block0_start_894_inst_ack_1 <= update_ack_unguarded(27);
      WPIPE_Block0_start_936_inst_ack_1 <= update_ack_unguarded(26);
      WPIPE_Block0_start_897_inst_ack_1 <= update_ack_unguarded(25);
      WPIPE_Block0_start_921_inst_ack_1 <= update_ack_unguarded(24);
      WPIPE_Block0_start_903_inst_ack_1 <= update_ack_unguarded(23);
      WPIPE_Block0_start_939_inst_ack_1 <= update_ack_unguarded(22);
      WPIPE_Block0_start_927_inst_ack_1 <= update_ack_unguarded(21);
      WPIPE_Block0_start_942_inst_ack_1 <= update_ack_unguarded(20);
      WPIPE_Block0_start_945_inst_ack_1 <= update_ack_unguarded(19);
      WPIPE_Block0_start_949_inst_ack_1 <= update_ack_unguarded(18);
      WPIPE_Block0_start_906_inst_ack_1 <= update_ack_unguarded(17);
      WPIPE_Block0_start_953_inst_ack_1 <= update_ack_unguarded(16);
      WPIPE_Block0_start_930_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Block0_start_957_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Block0_start_909_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_912_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_933_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_961_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_964_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_915_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_967_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_970_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_918_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_973_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_976_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_924_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_900_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_891_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      data_in <= call_35 & call92_258 & call10_73 & call46_173 & call19_98 & call106_267 & call55_198 & call101_264 & type_cast_947_wire_constant & type_cast_951_wire_constant & call14_85 & type_cast_955_wire_constant & call50_185 & type_cast_959_wire_constant & call28_123 & call23_110 & call97_261 & call115_283 & call110_270 & call37_148 & call124_308 & call119_295 & call32_135 & call133_333 & call128_320 & call41_160 & call5_60 & call2_48;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 8, num_reqs => 28, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_979_inst WPIPE_Block1_start_988_inst WPIPE_Block1_start_991_inst WPIPE_Block1_start_994_inst WPIPE_Block1_start_1000_inst WPIPE_Block1_start_997_inst WPIPE_Block1_start_1003_inst WPIPE_Block1_start_985_inst WPIPE_Block1_start_982_inst WPIPE_Block1_start_1006_inst WPIPE_Block1_start_1009_inst WPIPE_Block1_start_1012_inst WPIPE_Block1_start_1015_inst WPIPE_Block1_start_1018_inst WPIPE_Block1_start_1021_inst WPIPE_Block1_start_1024_inst WPIPE_Block1_start_1027_inst WPIPE_Block1_start_1030_inst WPIPE_Block1_start_1037_inst WPIPE_Block1_start_1050_inst WPIPE_Block1_start_1053_inst WPIPE_Block1_start_1056_inst WPIPE_Block1_start_1059_inst WPIPE_Block1_start_1062_inst WPIPE_Block1_start_1065_inst WPIPE_Block1_start_1068_inst WPIPE_Block1_start_1071_inst WPIPE_Block1_start_1074_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 27 downto 0);
      signal update_req, update_ack : BooleanArray( 27 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 27 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant inBUFs : IntegerArray(27 downto 0) := (27 => 0, 26 => 0, 25 => 0, 24 => 0, 23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      sample_req_unguarded(27) <= WPIPE_Block1_start_979_inst_req_0;
      sample_req_unguarded(26) <= WPIPE_Block1_start_988_inst_req_0;
      sample_req_unguarded(25) <= WPIPE_Block1_start_991_inst_req_0;
      sample_req_unguarded(24) <= WPIPE_Block1_start_994_inst_req_0;
      sample_req_unguarded(23) <= WPIPE_Block1_start_1000_inst_req_0;
      sample_req_unguarded(22) <= WPIPE_Block1_start_997_inst_req_0;
      sample_req_unguarded(21) <= WPIPE_Block1_start_1003_inst_req_0;
      sample_req_unguarded(20) <= WPIPE_Block1_start_985_inst_req_0;
      sample_req_unguarded(19) <= WPIPE_Block1_start_982_inst_req_0;
      sample_req_unguarded(18) <= WPIPE_Block1_start_1006_inst_req_0;
      sample_req_unguarded(17) <= WPIPE_Block1_start_1009_inst_req_0;
      sample_req_unguarded(16) <= WPIPE_Block1_start_1012_inst_req_0;
      sample_req_unguarded(15) <= WPIPE_Block1_start_1015_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Block1_start_1018_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Block1_start_1021_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1024_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1027_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1030_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1037_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1050_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1053_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1056_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1059_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1062_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1065_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1068_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1071_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1074_inst_req_0;
      WPIPE_Block1_start_979_inst_ack_0 <= sample_ack_unguarded(27);
      WPIPE_Block1_start_988_inst_ack_0 <= sample_ack_unguarded(26);
      WPIPE_Block1_start_991_inst_ack_0 <= sample_ack_unguarded(25);
      WPIPE_Block1_start_994_inst_ack_0 <= sample_ack_unguarded(24);
      WPIPE_Block1_start_1000_inst_ack_0 <= sample_ack_unguarded(23);
      WPIPE_Block1_start_997_inst_ack_0 <= sample_ack_unguarded(22);
      WPIPE_Block1_start_1003_inst_ack_0 <= sample_ack_unguarded(21);
      WPIPE_Block1_start_985_inst_ack_0 <= sample_ack_unguarded(20);
      WPIPE_Block1_start_982_inst_ack_0 <= sample_ack_unguarded(19);
      WPIPE_Block1_start_1006_inst_ack_0 <= sample_ack_unguarded(18);
      WPIPE_Block1_start_1009_inst_ack_0 <= sample_ack_unguarded(17);
      WPIPE_Block1_start_1012_inst_ack_0 <= sample_ack_unguarded(16);
      WPIPE_Block1_start_1015_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Block1_start_1018_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Block1_start_1021_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1024_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1027_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1030_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1037_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1050_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1053_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1056_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1059_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1062_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1065_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1068_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1071_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1074_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(27) <= WPIPE_Block1_start_979_inst_req_1;
      update_req_unguarded(26) <= WPIPE_Block1_start_988_inst_req_1;
      update_req_unguarded(25) <= WPIPE_Block1_start_991_inst_req_1;
      update_req_unguarded(24) <= WPIPE_Block1_start_994_inst_req_1;
      update_req_unguarded(23) <= WPIPE_Block1_start_1000_inst_req_1;
      update_req_unguarded(22) <= WPIPE_Block1_start_997_inst_req_1;
      update_req_unguarded(21) <= WPIPE_Block1_start_1003_inst_req_1;
      update_req_unguarded(20) <= WPIPE_Block1_start_985_inst_req_1;
      update_req_unguarded(19) <= WPIPE_Block1_start_982_inst_req_1;
      update_req_unguarded(18) <= WPIPE_Block1_start_1006_inst_req_1;
      update_req_unguarded(17) <= WPIPE_Block1_start_1009_inst_req_1;
      update_req_unguarded(16) <= WPIPE_Block1_start_1012_inst_req_1;
      update_req_unguarded(15) <= WPIPE_Block1_start_1015_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Block1_start_1018_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Block1_start_1021_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1024_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1027_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1030_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1037_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1050_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1053_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1056_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1059_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1062_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1065_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1068_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1071_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1074_inst_req_1;
      WPIPE_Block1_start_979_inst_ack_1 <= update_ack_unguarded(27);
      WPIPE_Block1_start_988_inst_ack_1 <= update_ack_unguarded(26);
      WPIPE_Block1_start_991_inst_ack_1 <= update_ack_unguarded(25);
      WPIPE_Block1_start_994_inst_ack_1 <= update_ack_unguarded(24);
      WPIPE_Block1_start_1000_inst_ack_1 <= update_ack_unguarded(23);
      WPIPE_Block1_start_997_inst_ack_1 <= update_ack_unguarded(22);
      WPIPE_Block1_start_1003_inst_ack_1 <= update_ack_unguarded(21);
      WPIPE_Block1_start_985_inst_ack_1 <= update_ack_unguarded(20);
      WPIPE_Block1_start_982_inst_ack_1 <= update_ack_unguarded(19);
      WPIPE_Block1_start_1006_inst_ack_1 <= update_ack_unguarded(18);
      WPIPE_Block1_start_1009_inst_ack_1 <= update_ack_unguarded(17);
      WPIPE_Block1_start_1012_inst_ack_1 <= update_ack_unguarded(16);
      WPIPE_Block1_start_1015_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Block1_start_1018_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Block1_start_1021_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1024_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1027_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1030_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1037_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1050_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1053_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1056_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1059_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1062_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1065_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1068_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1071_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1074_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      data_in <= call2_48 & call5_60 & call19_98 & call14_85 & call23_110 & call28_123 & call37_148 & call10_73 & call_35 & call32_135 & call46_173 & call41_160 & call55_198 & call50_185 & call97_261 & call92_258 & call106_267 & call101_264 & conv415_1036 & conv418_1049 & conv418_1049 & conv418_1049 & call115_283 & call110_270 & call124_308 & call119_295 & call133_333 & call128_320;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 8, num_reqs => 28, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1077_inst WPIPE_Block2_start_1080_inst WPIPE_Block2_start_1083_inst WPIPE_Block2_start_1086_inst WPIPE_Block2_start_1089_inst WPIPE_Block2_start_1092_inst WPIPE_Block2_start_1095_inst WPIPE_Block2_start_1098_inst WPIPE_Block2_start_1101_inst WPIPE_Block2_start_1104_inst WPIPE_Block2_start_1107_inst WPIPE_Block2_start_1110_inst WPIPE_Block2_start_1113_inst WPIPE_Block2_start_1116_inst WPIPE_Block2_start_1119_inst WPIPE_Block2_start_1122_inst WPIPE_Block2_start_1125_inst WPIPE_Block2_start_1128_inst WPIPE_Block2_start_1131_inst WPIPE_Block2_start_1145_inst WPIPE_Block2_start_1148_inst WPIPE_Block2_start_1151_inst WPIPE_Block2_start_1154_inst WPIPE_Block2_start_1157_inst WPIPE_Block2_start_1160_inst WPIPE_Block2_start_1163_inst WPIPE_Block2_start_1166_inst WPIPE_Block2_start_1169_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 27 downto 0);
      signal update_req, update_ack : BooleanArray( 27 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 27 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant inBUFs : IntegerArray(27 downto 0) := (27 => 0, 26 => 0, 25 => 0, 24 => 0, 23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      sample_req_unguarded(27) <= WPIPE_Block2_start_1077_inst_req_0;
      sample_req_unguarded(26) <= WPIPE_Block2_start_1080_inst_req_0;
      sample_req_unguarded(25) <= WPIPE_Block2_start_1083_inst_req_0;
      sample_req_unguarded(24) <= WPIPE_Block2_start_1086_inst_req_0;
      sample_req_unguarded(23) <= WPIPE_Block2_start_1089_inst_req_0;
      sample_req_unguarded(22) <= WPIPE_Block2_start_1092_inst_req_0;
      sample_req_unguarded(21) <= WPIPE_Block2_start_1095_inst_req_0;
      sample_req_unguarded(20) <= WPIPE_Block2_start_1098_inst_req_0;
      sample_req_unguarded(19) <= WPIPE_Block2_start_1101_inst_req_0;
      sample_req_unguarded(18) <= WPIPE_Block2_start_1104_inst_req_0;
      sample_req_unguarded(17) <= WPIPE_Block2_start_1107_inst_req_0;
      sample_req_unguarded(16) <= WPIPE_Block2_start_1110_inst_req_0;
      sample_req_unguarded(15) <= WPIPE_Block2_start_1113_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Block2_start_1116_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Block2_start_1119_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1122_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1125_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1128_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1131_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1145_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1148_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1151_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1154_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1157_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1160_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1163_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1166_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1169_inst_req_0;
      WPIPE_Block2_start_1077_inst_ack_0 <= sample_ack_unguarded(27);
      WPIPE_Block2_start_1080_inst_ack_0 <= sample_ack_unguarded(26);
      WPIPE_Block2_start_1083_inst_ack_0 <= sample_ack_unguarded(25);
      WPIPE_Block2_start_1086_inst_ack_0 <= sample_ack_unguarded(24);
      WPIPE_Block2_start_1089_inst_ack_0 <= sample_ack_unguarded(23);
      WPIPE_Block2_start_1092_inst_ack_0 <= sample_ack_unguarded(22);
      WPIPE_Block2_start_1095_inst_ack_0 <= sample_ack_unguarded(21);
      WPIPE_Block2_start_1098_inst_ack_0 <= sample_ack_unguarded(20);
      WPIPE_Block2_start_1101_inst_ack_0 <= sample_ack_unguarded(19);
      WPIPE_Block2_start_1104_inst_ack_0 <= sample_ack_unguarded(18);
      WPIPE_Block2_start_1107_inst_ack_0 <= sample_ack_unguarded(17);
      WPIPE_Block2_start_1110_inst_ack_0 <= sample_ack_unguarded(16);
      WPIPE_Block2_start_1113_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Block2_start_1116_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Block2_start_1119_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1122_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1125_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1128_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1131_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1145_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1148_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1151_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1154_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1157_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1160_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1163_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1166_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1169_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(27) <= WPIPE_Block2_start_1077_inst_req_1;
      update_req_unguarded(26) <= WPIPE_Block2_start_1080_inst_req_1;
      update_req_unguarded(25) <= WPIPE_Block2_start_1083_inst_req_1;
      update_req_unguarded(24) <= WPIPE_Block2_start_1086_inst_req_1;
      update_req_unguarded(23) <= WPIPE_Block2_start_1089_inst_req_1;
      update_req_unguarded(22) <= WPIPE_Block2_start_1092_inst_req_1;
      update_req_unguarded(21) <= WPIPE_Block2_start_1095_inst_req_1;
      update_req_unguarded(20) <= WPIPE_Block2_start_1098_inst_req_1;
      update_req_unguarded(19) <= WPIPE_Block2_start_1101_inst_req_1;
      update_req_unguarded(18) <= WPIPE_Block2_start_1104_inst_req_1;
      update_req_unguarded(17) <= WPIPE_Block2_start_1107_inst_req_1;
      update_req_unguarded(16) <= WPIPE_Block2_start_1110_inst_req_1;
      update_req_unguarded(15) <= WPIPE_Block2_start_1113_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Block2_start_1116_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Block2_start_1119_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1122_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1125_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1128_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1131_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1145_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1148_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1151_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1154_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1157_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1160_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1163_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1166_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1169_inst_req_1;
      WPIPE_Block2_start_1077_inst_ack_1 <= update_ack_unguarded(27);
      WPIPE_Block2_start_1080_inst_ack_1 <= update_ack_unguarded(26);
      WPIPE_Block2_start_1083_inst_ack_1 <= update_ack_unguarded(25);
      WPIPE_Block2_start_1086_inst_ack_1 <= update_ack_unguarded(24);
      WPIPE_Block2_start_1089_inst_ack_1 <= update_ack_unguarded(23);
      WPIPE_Block2_start_1092_inst_ack_1 <= update_ack_unguarded(22);
      WPIPE_Block2_start_1095_inst_ack_1 <= update_ack_unguarded(21);
      WPIPE_Block2_start_1098_inst_ack_1 <= update_ack_unguarded(20);
      WPIPE_Block2_start_1101_inst_ack_1 <= update_ack_unguarded(19);
      WPIPE_Block2_start_1104_inst_ack_1 <= update_ack_unguarded(18);
      WPIPE_Block2_start_1107_inst_ack_1 <= update_ack_unguarded(17);
      WPIPE_Block2_start_1110_inst_ack_1 <= update_ack_unguarded(16);
      WPIPE_Block2_start_1113_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Block2_start_1116_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Block2_start_1119_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1122_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1125_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1128_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1131_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1145_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1148_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1151_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1154_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1157_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1160_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1163_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1166_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1169_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      data_in <= call2_48 & call_35 & call10_73 & call5_60 & call19_98 & call14_85 & call28_123 & call23_110 & call37_148 & call32_135 & call46_173 & call41_160 & call55_198 & call50_185 & call97_261 & call92_258 & call106_267 & call101_264 & type_cast_1133_wire_constant & conv501_1144 & conv501_1144 & conv501_1144 & call115_283 & call110_270 & call124_308 & call119_295 & call133_333 & call128_320;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 8, num_reqs => 28, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1172_inst WPIPE_Block3_start_1175_inst WPIPE_Block3_start_1178_inst WPIPE_Block3_start_1181_inst WPIPE_Block3_start_1184_inst WPIPE_Block3_start_1187_inst WPIPE_Block3_start_1190_inst WPIPE_Block3_start_1193_inst WPIPE_Block3_start_1196_inst WPIPE_Block3_start_1199_inst WPIPE_Block3_start_1202_inst WPIPE_Block3_start_1205_inst WPIPE_Block3_start_1208_inst WPIPE_Block3_start_1211_inst WPIPE_Block3_start_1214_inst WPIPE_Block3_start_1217_inst WPIPE_Block3_start_1220_inst WPIPE_Block3_start_1223_inst WPIPE_Block3_start_1226_inst WPIPE_Block3_start_1240_inst WPIPE_Block3_start_1243_inst WPIPE_Block3_start_1246_inst WPIPE_Block3_start_1249_inst WPIPE_Block3_start_1252_inst WPIPE_Block3_start_1255_inst WPIPE_Block3_start_1258_inst WPIPE_Block3_start_1261_inst WPIPE_Block3_start_1264_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 27 downto 0);
      signal update_req, update_ack : BooleanArray( 27 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 27 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant inBUFs : IntegerArray(27 downto 0) := (27 => 0, 26 => 0, 25 => 0, 24 => 0, 23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      sample_req_unguarded(27) <= WPIPE_Block3_start_1172_inst_req_0;
      sample_req_unguarded(26) <= WPIPE_Block3_start_1175_inst_req_0;
      sample_req_unguarded(25) <= WPIPE_Block3_start_1178_inst_req_0;
      sample_req_unguarded(24) <= WPIPE_Block3_start_1181_inst_req_0;
      sample_req_unguarded(23) <= WPIPE_Block3_start_1184_inst_req_0;
      sample_req_unguarded(22) <= WPIPE_Block3_start_1187_inst_req_0;
      sample_req_unguarded(21) <= WPIPE_Block3_start_1190_inst_req_0;
      sample_req_unguarded(20) <= WPIPE_Block3_start_1193_inst_req_0;
      sample_req_unguarded(19) <= WPIPE_Block3_start_1196_inst_req_0;
      sample_req_unguarded(18) <= WPIPE_Block3_start_1199_inst_req_0;
      sample_req_unguarded(17) <= WPIPE_Block3_start_1202_inst_req_0;
      sample_req_unguarded(16) <= WPIPE_Block3_start_1205_inst_req_0;
      sample_req_unguarded(15) <= WPIPE_Block3_start_1208_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Block3_start_1211_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Block3_start_1214_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1217_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1220_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1223_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1226_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1240_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1243_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1246_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1249_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1252_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1255_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1258_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1261_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1264_inst_req_0;
      WPIPE_Block3_start_1172_inst_ack_0 <= sample_ack_unguarded(27);
      WPIPE_Block3_start_1175_inst_ack_0 <= sample_ack_unguarded(26);
      WPIPE_Block3_start_1178_inst_ack_0 <= sample_ack_unguarded(25);
      WPIPE_Block3_start_1181_inst_ack_0 <= sample_ack_unguarded(24);
      WPIPE_Block3_start_1184_inst_ack_0 <= sample_ack_unguarded(23);
      WPIPE_Block3_start_1187_inst_ack_0 <= sample_ack_unguarded(22);
      WPIPE_Block3_start_1190_inst_ack_0 <= sample_ack_unguarded(21);
      WPIPE_Block3_start_1193_inst_ack_0 <= sample_ack_unguarded(20);
      WPIPE_Block3_start_1196_inst_ack_0 <= sample_ack_unguarded(19);
      WPIPE_Block3_start_1199_inst_ack_0 <= sample_ack_unguarded(18);
      WPIPE_Block3_start_1202_inst_ack_0 <= sample_ack_unguarded(17);
      WPIPE_Block3_start_1205_inst_ack_0 <= sample_ack_unguarded(16);
      WPIPE_Block3_start_1208_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Block3_start_1211_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Block3_start_1214_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1217_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1220_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1223_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1226_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1240_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1243_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1246_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1249_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1252_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1255_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1258_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1261_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1264_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(27) <= WPIPE_Block3_start_1172_inst_req_1;
      update_req_unguarded(26) <= WPIPE_Block3_start_1175_inst_req_1;
      update_req_unguarded(25) <= WPIPE_Block3_start_1178_inst_req_1;
      update_req_unguarded(24) <= WPIPE_Block3_start_1181_inst_req_1;
      update_req_unguarded(23) <= WPIPE_Block3_start_1184_inst_req_1;
      update_req_unguarded(22) <= WPIPE_Block3_start_1187_inst_req_1;
      update_req_unguarded(21) <= WPIPE_Block3_start_1190_inst_req_1;
      update_req_unguarded(20) <= WPIPE_Block3_start_1193_inst_req_1;
      update_req_unguarded(19) <= WPIPE_Block3_start_1196_inst_req_1;
      update_req_unguarded(18) <= WPIPE_Block3_start_1199_inst_req_1;
      update_req_unguarded(17) <= WPIPE_Block3_start_1202_inst_req_1;
      update_req_unguarded(16) <= WPIPE_Block3_start_1205_inst_req_1;
      update_req_unguarded(15) <= WPIPE_Block3_start_1208_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Block3_start_1211_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Block3_start_1214_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1217_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1220_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1223_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1226_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1240_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1243_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1246_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1249_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1252_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1255_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1258_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1261_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1264_inst_req_1;
      WPIPE_Block3_start_1172_inst_ack_1 <= update_ack_unguarded(27);
      WPIPE_Block3_start_1175_inst_ack_1 <= update_ack_unguarded(26);
      WPIPE_Block3_start_1178_inst_ack_1 <= update_ack_unguarded(25);
      WPIPE_Block3_start_1181_inst_ack_1 <= update_ack_unguarded(24);
      WPIPE_Block3_start_1184_inst_ack_1 <= update_ack_unguarded(23);
      WPIPE_Block3_start_1187_inst_ack_1 <= update_ack_unguarded(22);
      WPIPE_Block3_start_1190_inst_ack_1 <= update_ack_unguarded(21);
      WPIPE_Block3_start_1193_inst_ack_1 <= update_ack_unguarded(20);
      WPIPE_Block3_start_1196_inst_ack_1 <= update_ack_unguarded(19);
      WPIPE_Block3_start_1199_inst_ack_1 <= update_ack_unguarded(18);
      WPIPE_Block3_start_1202_inst_ack_1 <= update_ack_unguarded(17);
      WPIPE_Block3_start_1205_inst_ack_1 <= update_ack_unguarded(16);
      WPIPE_Block3_start_1208_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Block3_start_1211_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Block3_start_1214_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1217_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1220_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1223_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1226_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1240_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1243_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1246_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1249_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1252_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1255_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1258_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1261_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1264_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      data_in <= call2_48 & call_35 & call10_73 & call5_60 & call19_98 & call14_85 & call28_123 & call23_110 & call37_148 & call32_135 & call46_173 & call41_160 & call55_198 & call50_185 & call97_261 & call92_258 & call106_267 & call101_264 & type_cast_1228_wire_constant & conv584_1239 & conv584_1239 & conv584_1239 & call115_283 & call110_270 & call124_308 & call119_295 & call133_333 & call128_320;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 8, num_reqs => 28, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1433_inst WPIPE_ConvTranspose_output_pipe_1436_inst WPIPE_ConvTranspose_output_pipe_1439_inst WPIPE_ConvTranspose_output_pipe_1442_inst WPIPE_ConvTranspose_output_pipe_1445_inst WPIPE_ConvTranspose_output_pipe_1448_inst WPIPE_ConvTranspose_output_pipe_1451_inst WPIPE_ConvTranspose_output_pipe_1454_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1433_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1436_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1439_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1442_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1445_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1448_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1451_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1454_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1433_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1436_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1439_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1442_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1445_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1433_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1436_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1439_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1442_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1445_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1448_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1451_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1454_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1433_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1436_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1439_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1442_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1445_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv681_1432 & conv675_1422 & conv669_1412 & conv663_1402 & conv657_1392 & conv651_1382 & conv645_1372 & conv639_1362;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_elapsed_time_pipe_1292_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1292_inst_req_0;
      WPIPE_elapsed_time_pipe_1292_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1292_inst_req_1;
      WPIPE_elapsed_time_pipe_1292_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1291;
      elapsed_time_pipe_write_5_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_5: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared call operator group (0) : call_stmt_884_call call_stmt_1281_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_884_call_req_0;
      reqL_unguarded(0) <= call_stmt_1281_call_req_0;
      call_stmt_884_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1281_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_884_call_req_1;
      reqR_unguarded(0) <= call_stmt_1281_call_req_1;
      call_stmt_884_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1281_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call275_884 <= data_out(127 downto 64);
      call618_1281 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_4108_start: Boolean;
  signal convTransposeA_CP_4108_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1551_inst_ack_1 : boolean;
  signal type_cast_1570_inst_req_1 : boolean;
  signal type_cast_1551_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1604_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1604_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1622_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1604_inst_req_0 : boolean;
  signal type_cast_1551_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1579_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1604_inst_req_1 : boolean;
  signal type_cast_1595_inst_ack_1 : boolean;
  signal type_cast_1639_inst_ack_0 : boolean;
  signal type_cast_1570_inst_ack_0 : boolean;
  signal type_cast_1570_inst_ack_1 : boolean;
  signal type_cast_1595_inst_req_1 : boolean;
  signal type_cast_1570_inst_req_0 : boolean;
  signal type_cast_1551_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1559_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1562_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1562_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1647_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1562_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1635_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1635_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1579_inst_ack_1 : boolean;
  signal type_cast_1608_inst_ack_0 : boolean;
  signal type_cast_1608_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1579_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1562_inst_ack_1 : boolean;
  signal type_cast_1651_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1559_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1559_inst_ack_1 : boolean;
  signal type_cast_1664_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1579_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1672_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1647_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1622_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1660_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1559_inst_ack_0 : boolean;
  signal type_cast_1608_inst_req_1 : boolean;
  signal type_cast_1608_inst_ack_1 : boolean;
  signal type_cast_1595_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1622_inst_ack_0 : boolean;
  signal type_cast_1595_inst_req_0 : boolean;
  signal type_cast_1664_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1622_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1635_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1685_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1635_inst_req_0 : boolean;
  signal type_cast_1664_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1685_inst_req_0 : boolean;
  signal type_cast_1651_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1565_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1685_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1565_inst_req_1 : boolean;
  signal type_cast_1583_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1565_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1616_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1616_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1565_inst_req_0 : boolean;
  signal type_cast_1639_inst_ack_1 : boolean;
  signal type_cast_1488_inst_req_0 : boolean;
  signal type_cast_1488_inst_ack_0 : boolean;
  signal type_cast_1488_inst_req_1 : boolean;
  signal type_cast_1488_inst_ack_1 : boolean;
  signal type_cast_1689_inst_req_0 : boolean;
  signal type_cast_1689_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1660_inst_ack_0 : boolean;
  signal type_cast_1583_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1672_inst_req_0 : boolean;
  signal type_cast_1651_inst_ack_0 : boolean;
  signal type_cast_1676_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1660_inst_req_1 : boolean;
  signal type_cast_1639_inst_req_0 : boolean;
  signal type_cast_1676_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1660_inst_ack_1 : boolean;
  signal type_cast_1583_inst_ack_0 : boolean;
  signal type_cast_1664_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1672_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1672_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1685_inst_ack_1 : boolean;
  signal type_cast_1651_inst_req_0 : boolean;
  signal type_cast_1676_inst_req_0 : boolean;
  signal type_cast_1676_inst_ack_0 : boolean;
  signal type_cast_1583_inst_req_1 : boolean;
  signal type_cast_1626_inst_ack_1 : boolean;
  signal type_cast_1626_inst_req_1 : boolean;
  signal type_cast_1626_inst_ack_0 : boolean;
  signal type_cast_1626_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1484_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1484_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1484_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1484_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1497_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1497_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1497_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1497_inst_ack_1 : boolean;
  signal type_cast_1501_inst_req_0 : boolean;
  signal type_cast_1501_inst_ack_0 : boolean;
  signal type_cast_1501_inst_req_1 : boolean;
  signal type_cast_1501_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1509_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1509_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1509_inst_ack_1 : boolean;
  signal type_cast_1513_inst_req_0 : boolean;
  signal type_cast_1513_inst_ack_0 : boolean;
  signal type_cast_1513_inst_req_1 : boolean;
  signal type_cast_1513_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1647_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1619_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1591_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1619_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1591_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1522_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1522_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1522_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1522_inst_ack_1 : boolean;
  signal type_cast_1639_inst_req_1 : boolean;
  signal type_cast_1526_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1616_inst_ack_0 : boolean;
  signal type_cast_1526_inst_ack_0 : boolean;
  signal type_cast_1526_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1616_inst_req_0 : boolean;
  signal type_cast_1526_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1547_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1647_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1619_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1619_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1591_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1591_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1534_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1534_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1547_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1534_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1534_inst_ack_1 : boolean;
  signal type_cast_1538_inst_req_0 : boolean;
  signal type_cast_1538_inst_ack_0 : boolean;
  signal type_cast_1538_inst_req_1 : boolean;
  signal type_cast_1538_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1547_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1547_inst_ack_0 : boolean;
  signal type_cast_1689_inst_req_1 : boolean;
  signal type_cast_1689_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1703_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1703_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1703_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1703_inst_ack_1 : boolean;
  signal type_cast_1707_inst_req_0 : boolean;
  signal type_cast_1707_inst_ack_0 : boolean;
  signal type_cast_1707_inst_req_1 : boolean;
  signal type_cast_1707_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1721_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1721_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1721_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1721_inst_ack_1 : boolean;
  signal type_cast_1725_inst_req_0 : boolean;
  signal type_cast_1725_inst_ack_0 : boolean;
  signal type_cast_1725_inst_req_1 : boolean;
  signal type_cast_1725_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1733_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1733_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1733_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1733_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1736_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1736_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1736_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1736_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1739_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1739_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1739_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1739_inst_ack_1 : boolean;
  signal type_cast_1743_inst_req_0 : boolean;
  signal type_cast_1743_inst_ack_0 : boolean;
  signal type_cast_1743_inst_req_1 : boolean;
  signal type_cast_1743_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1752_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1752_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1752_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1752_inst_ack_1 : boolean;
  signal type_cast_1756_inst_req_0 : boolean;
  signal type_cast_1756_inst_ack_0 : boolean;
  signal type_cast_1756_inst_req_1 : boolean;
  signal type_cast_1756_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1764_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1764_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1764_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1764_inst_ack_1 : boolean;
  signal type_cast_1768_inst_req_0 : boolean;
  signal type_cast_1768_inst_ack_0 : boolean;
  signal type_cast_1768_inst_req_1 : boolean;
  signal type_cast_1768_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1777_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1777_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1777_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1777_inst_ack_1 : boolean;
  signal type_cast_1781_inst_req_0 : boolean;
  signal type_cast_1781_inst_ack_0 : boolean;
  signal type_cast_1781_inst_req_1 : boolean;
  signal type_cast_1781_inst_ack_1 : boolean;
  signal type_cast_1881_inst_req_0 : boolean;
  signal type_cast_1881_inst_ack_0 : boolean;
  signal type_cast_1881_inst_req_1 : boolean;
  signal type_cast_1881_inst_ack_1 : boolean;
  signal type_cast_1885_inst_req_0 : boolean;
  signal type_cast_1885_inst_ack_0 : boolean;
  signal type_cast_1885_inst_req_1 : boolean;
  signal type_cast_1885_inst_ack_1 : boolean;
  signal phi_stmt_2045_req_1 : boolean;
  signal type_cast_1889_inst_req_0 : boolean;
  signal type_cast_1889_inst_ack_0 : boolean;
  signal type_cast_1889_inst_req_1 : boolean;
  signal type_cast_1889_inst_ack_1 : boolean;
  signal type_cast_2050_inst_ack_1 : boolean;
  signal type_cast_1919_inst_req_0 : boolean;
  signal type_cast_1919_inst_ack_0 : boolean;
  signal type_cast_1919_inst_req_1 : boolean;
  signal type_cast_1919_inst_ack_1 : boolean;
  signal type_cast_2050_inst_req_1 : boolean;
  signal type_cast_2050_inst_ack_0 : boolean;
  signal type_cast_2050_inst_req_0 : boolean;
  signal array_obj_ref_1925_index_offset_req_0 : boolean;
  signal array_obj_ref_1925_index_offset_ack_0 : boolean;
  signal phi_stmt_2045_req_0 : boolean;
  signal array_obj_ref_1925_index_offset_req_1 : boolean;
  signal array_obj_ref_1925_index_offset_ack_1 : boolean;
  signal type_cast_2048_inst_ack_1 : boolean;
  signal addr_of_1926_final_reg_req_0 : boolean;
  signal addr_of_1926_final_reg_ack_0 : boolean;
  signal addr_of_1926_final_reg_req_1 : boolean;
  signal addr_of_1926_final_reg_ack_1 : boolean;
  signal type_cast_2044_inst_ack_0 : boolean;
  signal type_cast_2044_inst_req_0 : boolean;
  signal ptr_deref_1930_load_0_req_0 : boolean;
  signal ptr_deref_1930_load_0_ack_0 : boolean;
  signal type_cast_2048_inst_req_0 : boolean;
  signal ptr_deref_1930_load_0_req_1 : boolean;
  signal ptr_deref_1930_load_0_ack_1 : boolean;
  signal array_obj_ref_1948_index_offset_req_0 : boolean;
  signal array_obj_ref_1948_index_offset_ack_0 : boolean;
  signal type_cast_2048_inst_req_1 : boolean;
  signal array_obj_ref_1948_index_offset_req_1 : boolean;
  signal array_obj_ref_1948_index_offset_ack_1 : boolean;
  signal addr_of_1949_final_reg_req_0 : boolean;
  signal phi_stmt_2045_ack_0 : boolean;
  signal addr_of_1949_final_reg_ack_0 : boolean;
  signal addr_of_1949_final_reg_req_1 : boolean;
  signal phi_stmt_2039_ack_0 : boolean;
  signal addr_of_1949_final_reg_ack_1 : boolean;
  signal phi_stmt_2032_ack_0 : boolean;
  signal phi_stmt_2032_req_1 : boolean;
  signal phi_stmt_2039_req_0 : boolean;
  signal phi_stmt_2032_req_0 : boolean;
  signal ptr_deref_1952_store_0_req_0 : boolean;
  signal ptr_deref_1952_store_0_ack_0 : boolean;
  signal type_cast_2042_inst_ack_1 : boolean;
  signal ptr_deref_1952_store_0_req_1 : boolean;
  signal ptr_deref_1952_store_0_ack_1 : boolean;
  signal type_cast_1957_inst_req_0 : boolean;
  signal type_cast_2035_inst_ack_1 : boolean;
  signal type_cast_1957_inst_ack_0 : boolean;
  signal type_cast_1957_inst_req_1 : boolean;
  signal type_cast_2035_inst_req_1 : boolean;
  signal type_cast_1957_inst_ack_1 : boolean;
  signal type_cast_2042_inst_req_1 : boolean;
  signal if_stmt_1970_branch_req_0 : boolean;
  signal phi_stmt_2039_req_1 : boolean;
  signal if_stmt_1970_branch_ack_1 : boolean;
  signal if_stmt_1970_branch_ack_0 : boolean;
  signal type_cast_2042_inst_ack_0 : boolean;
  signal type_cast_2042_inst_req_0 : boolean;
  signal type_cast_1993_inst_req_0 : boolean;
  signal type_cast_1993_inst_ack_0 : boolean;
  signal type_cast_1993_inst_req_1 : boolean;
  signal type_cast_1993_inst_ack_1 : boolean;
  signal type_cast_2044_inst_ack_1 : boolean;
  signal type_cast_2002_inst_req_0 : boolean;
  signal type_cast_2035_inst_ack_0 : boolean;
  signal type_cast_2002_inst_ack_0 : boolean;
  signal type_cast_2002_inst_req_1 : boolean;
  signal type_cast_2035_inst_req_0 : boolean;
  signal type_cast_2002_inst_ack_1 : boolean;
  signal type_cast_2044_inst_req_1 : boolean;
  signal type_cast_2018_inst_req_0 : boolean;
  signal type_cast_2018_inst_ack_0 : boolean;
  signal type_cast_2018_inst_req_1 : boolean;
  signal type_cast_2018_inst_ack_1 : boolean;
  signal type_cast_2048_inst_ack_0 : boolean;
  signal if_stmt_2025_branch_req_0 : boolean;
  signal if_stmt_2025_branch_ack_1 : boolean;
  signal if_stmt_2025_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_2061_inst_req_0 : boolean;
  signal WPIPE_Block0_done_2061_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_2061_inst_req_1 : boolean;
  signal WPIPE_Block0_done_2061_inst_ack_1 : boolean;
  signal phi_stmt_1819_req_0 : boolean;
  signal phi_stmt_1826_req_0 : boolean;
  signal phi_stmt_1833_req_0 : boolean;
  signal phi_stmt_1840_req_0 : boolean;
  signal type_cast_1825_inst_req_0 : boolean;
  signal type_cast_1825_inst_ack_0 : boolean;
  signal type_cast_1825_inst_req_1 : boolean;
  signal type_cast_1825_inst_ack_1 : boolean;
  signal phi_stmt_1819_req_1 : boolean;
  signal type_cast_1832_inst_req_0 : boolean;
  signal type_cast_1832_inst_ack_0 : boolean;
  signal type_cast_1832_inst_req_1 : boolean;
  signal type_cast_1832_inst_ack_1 : boolean;
  signal phi_stmt_1826_req_1 : boolean;
  signal type_cast_1839_inst_req_0 : boolean;
  signal type_cast_1839_inst_ack_0 : boolean;
  signal type_cast_1839_inst_req_1 : boolean;
  signal type_cast_1839_inst_ack_1 : boolean;
  signal phi_stmt_1833_req_1 : boolean;
  signal type_cast_1846_inst_req_0 : boolean;
  signal type_cast_1846_inst_ack_0 : boolean;
  signal type_cast_1846_inst_req_1 : boolean;
  signal type_cast_1846_inst_ack_1 : boolean;
  signal phi_stmt_1840_req_1 : boolean;
  signal phi_stmt_1819_ack_0 : boolean;
  signal phi_stmt_1826_ack_0 : boolean;
  signal phi_stmt_1833_ack_0 : boolean;
  signal phi_stmt_1840_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_4108_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_4108_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_4108_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_4108_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_4108: Block -- control-path 
    signal convTransposeA_CP_4108_elements: BooleanArray(186 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_4108_elements(0) <= convTransposeA_CP_4108_start;
    convTransposeA_CP_4108_symbol <= convTransposeA_CP_4108_elements(139);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	41 
    -- CP-element group 0:  members (74) 
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1482/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/branch_block_stmt_1482__entry__
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787__entry__
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_Update/cr
      -- 
    cr_4371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1570_inst_req_1); -- 
    cr_4315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1551_inst_req_1); -- 
    cr_4427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1595_inst_req_1); -- 
    cr_4455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1608_inst_req_1); -- 
    cr_4595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1664_inst_req_1); -- 
    cr_4567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1651_inst_req_1); -- 
    cr_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1488_inst_req_1); -- 
    cr_4623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1676_inst_req_1); -- 
    cr_4399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1583_inst_req_1); -- 
    cr_4511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1626_inst_req_1); -- 
    rr_4156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => RPIPE_Block0_start_1484_inst_req_0); -- 
    cr_4203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1501_inst_req_1); -- 
    cr_4231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1513_inst_req_1); -- 
    cr_4539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1639_inst_req_1); -- 
    cr_4259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1526_inst_req_1); -- 
    cr_4287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1538_inst_req_1); -- 
    cr_4651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1689_inst_req_1); -- 
    cr_4679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1707_inst_req_1); -- 
    cr_4707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1725_inst_req_1); -- 
    cr_4763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1743_inst_req_1); -- 
    cr_4791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1756_inst_req_1); -- 
    cr_4819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1768_inst_req_1); -- 
    cr_4847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(0), ack => type_cast_1781_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	186 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	145 
    -- CP-element group 1: 	146 
    -- CP-element group 1: 	148 
    -- CP-element group 1: 	149 
    -- CP-element group 1: 	151 
    -- CP-element group 1: 	152 
    -- CP-element group 1: 	154 
    -- CP-element group 1: 	155 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1482/merge_stmt_2031__exit__
      -- CP-element group 1: 	 branch_block_stmt_1482/assign_stmt_2057__entry__
      -- CP-element group 1: 	 branch_block_stmt_1482/assign_stmt_2057__exit__
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1482/assign_stmt_2057/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/assign_stmt_2057/$exit
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/Update/cr
      -- 
    rr_5276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(1), ack => type_cast_1825_inst_req_0); -- 
    cr_5281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(1), ack => type_cast_1825_inst_req_1); -- 
    rr_5299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(1), ack => type_cast_1832_inst_req_0); -- 
    cr_5304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(1), ack => type_cast_1832_inst_req_1); -- 
    rr_5322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(1), ack => type_cast_1839_inst_req_0); -- 
    cr_5327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(1), ack => type_cast_1839_inst_req_1); -- 
    rr_5345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(1), ack => type_cast_1846_inst_req_0); -- 
    cr_5350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(1), ack => type_cast_1846_inst_req_1); -- 
    convTransposeA_CP_4108_elements(1) <= convTransposeA_CP_4108_elements(186);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_Update/cr
      -- 
    ra_4157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1484_inst_ack_0, ack => convTransposeA_CP_4108_elements(2)); -- 
    cr_4161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(2), ack => RPIPE_Block0_start_1484_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1484_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_Sample/rr
      -- 
    ca_4162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1484_inst_ack_1, ack => convTransposeA_CP_4108_elements(3)); -- 
    rr_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(3), ack => type_cast_1488_inst_req_0); -- 
    rr_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(3), ack => RPIPE_Block0_start_1497_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_sample_completed_
      -- 
    ra_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_0, ack => convTransposeA_CP_4108_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	102 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1488_update_completed_
      -- 
    ca_4176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1488_inst_ack_1, ack => convTransposeA_CP_4108_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_Update/cr
      -- 
    ra_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1497_inst_ack_0, ack => convTransposeA_CP_4108_elements(6)); -- 
    cr_4189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(6), ack => RPIPE_Block0_start_1497_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1497_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_Sample/rr
      -- 
    ca_4190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1497_inst_ack_1, ack => convTransposeA_CP_4108_elements(7)); -- 
    rr_4198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(7), ack => type_cast_1501_inst_req_0); -- 
    rr_4212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(7), ack => RPIPE_Block0_start_1509_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_Sample/ra
      -- 
    ra_4199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1501_inst_ack_0, ack => convTransposeA_CP_4108_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	102 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1501_Update/ca
      -- 
    ca_4204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1501_inst_ack_1, ack => convTransposeA_CP_4108_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_Update/cr
      -- 
    ra_4213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1509_inst_ack_0, ack => convTransposeA_CP_4108_elements(10)); -- 
    cr_4217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(10), ack => RPIPE_Block0_start_1509_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1509_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_Sample/rr
      -- 
    ca_4218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1509_inst_ack_1, ack => convTransposeA_CP_4108_elements(11)); -- 
    rr_4226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(11), ack => type_cast_1513_inst_req_0); -- 
    rr_4240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(11), ack => RPIPE_Block0_start_1522_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_Sample/ra
      -- 
    ra_4227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1513_inst_ack_0, ack => convTransposeA_CP_4108_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	102 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1513_Update/ca
      -- 
    ca_4232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1513_inst_ack_1, ack => convTransposeA_CP_4108_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_Update/cr
      -- 
    ra_4241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1522_inst_ack_0, ack => convTransposeA_CP_4108_elements(14)); -- 
    cr_4245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(14), ack => RPIPE_Block0_start_1522_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1522_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_Sample/rr
      -- 
    ca_4246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1522_inst_ack_1, ack => convTransposeA_CP_4108_elements(15)); -- 
    rr_4254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(15), ack => type_cast_1526_inst_req_0); -- 
    rr_4268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(15), ack => RPIPE_Block0_start_1534_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_Sample/ra
      -- 
    ra_4255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1526_inst_ack_0, ack => convTransposeA_CP_4108_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	102 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1526_Update/ca
      -- 
    ca_4260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1526_inst_ack_1, ack => convTransposeA_CP_4108_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_Update/cr
      -- 
    ra_4269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1534_inst_ack_0, ack => convTransposeA_CP_4108_elements(18)); -- 
    cr_4273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(18), ack => RPIPE_Block0_start_1534_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1534_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_Sample/rr
      -- 
    ca_4274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1534_inst_ack_1, ack => convTransposeA_CP_4108_elements(19)); -- 
    rr_4282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(19), ack => type_cast_1538_inst_req_0); -- 
    rr_4296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(19), ack => RPIPE_Block0_start_1547_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_Sample/ra
      -- 
    ra_4283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_0, ack => convTransposeA_CP_4108_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	102 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1538_Update/ca
      -- 
    ca_4288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1538_inst_ack_1, ack => convTransposeA_CP_4108_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_Sample/ra
      -- 
    ra_4297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1547_inst_ack_0, ack => convTransposeA_CP_4108_elements(22)); -- 
    cr_4301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(22), ack => RPIPE_Block0_start_1547_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1547_update_completed_
      -- 
    ca_4302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1547_inst_ack_1, ack => convTransposeA_CP_4108_elements(23)); -- 
    rr_4310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(23), ack => type_cast_1551_inst_req_0); -- 
    rr_4324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(23), ack => RPIPE_Block0_start_1559_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_sample_completed_
      -- 
    ra_4311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1551_inst_ack_0, ack => convTransposeA_CP_4108_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	102 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1551_update_completed_
      -- 
    ca_4316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1551_inst_ack_1, ack => convTransposeA_CP_4108_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_update_start_
      -- 
    ra_4325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1559_inst_ack_0, ack => convTransposeA_CP_4108_elements(26)); -- 
    cr_4329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(26), ack => RPIPE_Block0_start_1559_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1559_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_sample_start_
      -- 
    ca_4330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1559_inst_ack_1, ack => convTransposeA_CP_4108_elements(27)); -- 
    rr_4338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(27), ack => RPIPE_Block0_start_1562_inst_req_0); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_update_start_
      -- 
    ra_4339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1562_inst_ack_0, ack => convTransposeA_CP_4108_elements(28)); -- 
    cr_4343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(28), ack => RPIPE_Block0_start_1562_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1562_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_Sample/$entry
      -- 
    ca_4344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1562_inst_ack_1, ack => convTransposeA_CP_4108_elements(29)); -- 
    rr_4352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(29), ack => RPIPE_Block0_start_1565_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_update_start_
      -- 
    ra_4353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1565_inst_ack_0, ack => convTransposeA_CP_4108_elements(30)); -- 
    cr_4357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(30), ack => RPIPE_Block0_start_1565_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1565_update_completed_
      -- 
    ca_4358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1565_inst_ack_1, ack => convTransposeA_CP_4108_elements(31)); -- 
    rr_4366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(31), ack => type_cast_1570_inst_req_0); -- 
    rr_4380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(31), ack => RPIPE_Block0_start_1579_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_sample_completed_
      -- 
    ra_4367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_0, ack => convTransposeA_CP_4108_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	102 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1570_update_completed_
      -- 
    ca_4372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_1, ack => convTransposeA_CP_4108_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_Update/$entry
      -- 
    ra_4381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1579_inst_ack_0, ack => convTransposeA_CP_4108_elements(34)); -- 
    cr_4385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(34), ack => RPIPE_Block0_start_1579_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1579_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_Sample/rr
      -- 
    ca_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1579_inst_ack_1, ack => convTransposeA_CP_4108_elements(35)); -- 
    rr_4394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(35), ack => type_cast_1583_inst_req_0); -- 
    rr_4408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(35), ack => RPIPE_Block0_start_1591_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_Sample/ra
      -- 
    ra_4395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1583_inst_ack_0, ack => convTransposeA_CP_4108_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	102 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1583_Update/ca
      -- 
    ca_4400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1583_inst_ack_1, ack => convTransposeA_CP_4108_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_Sample/$exit
      -- 
    ra_4409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1591_inst_ack_0, ack => convTransposeA_CP_4108_elements(38)); -- 
    cr_4413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(38), ack => RPIPE_Block0_start_1591_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1591_Update/$exit
      -- 
    ca_4414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1591_inst_ack_1, ack => convTransposeA_CP_4108_elements(39)); -- 
    rr_4422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(39), ack => type_cast_1595_inst_req_0); -- 
    rr_4436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(39), ack => RPIPE_Block0_start_1604_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_Sample/ra
      -- CP-element group 40: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_sample_completed_
      -- 
    ra_4423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1595_inst_ack_0, ack => convTransposeA_CP_4108_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	102 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_Update/ca
      -- CP-element group 41: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1595_update_completed_
      -- 
    ca_4428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1595_inst_ack_1, ack => convTransposeA_CP_4108_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_update_start_
      -- CP-element group 42: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_Update/cr
      -- CP-element group 42: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_Sample/$exit
      -- 
    ra_4437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1604_inst_ack_0, ack => convTransposeA_CP_4108_elements(42)); -- 
    cr_4441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(42), ack => RPIPE_Block0_start_1604_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	46 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1604_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_Sample/rr
      -- 
    ca_4442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1604_inst_ack_1, ack => convTransposeA_CP_4108_elements(43)); -- 
    rr_4464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(43), ack => RPIPE_Block0_start_1616_inst_req_0); -- 
    rr_4450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(43), ack => type_cast_1608_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_Sample/$exit
      -- 
    ra_4451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1608_inst_ack_0, ack => convTransposeA_CP_4108_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	102 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1608_Update/ca
      -- 
    ca_4456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1608_inst_ack_1, ack => convTransposeA_CP_4108_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_Update/cr
      -- CP-element group 46: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_Sample/$exit
      -- 
    ra_4465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1616_inst_ack_0, ack => convTransposeA_CP_4108_elements(46)); -- 
    cr_4469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(46), ack => RPIPE_Block0_start_1616_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1616_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_Sample/rr
      -- 
    ca_4470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1616_inst_ack_1, ack => convTransposeA_CP_4108_elements(47)); -- 
    rr_4478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(47), ack => RPIPE_Block0_start_1619_inst_req_0); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_Update/cr
      -- CP-element group 48: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_Sample/ra
      -- 
    ra_4479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1619_inst_ack_0, ack => convTransposeA_CP_4108_elements(48)); -- 
    cr_4483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(48), ack => RPIPE_Block0_start_1619_inst_req_1); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1619_Update/$exit
      -- 
    ca_4484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1619_inst_ack_1, ack => convTransposeA_CP_4108_elements(49)); -- 
    rr_4492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(49), ack => RPIPE_Block0_start_1622_inst_req_0); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_Update/cr
      -- CP-element group 50: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_sample_completed_
      -- 
    ra_4493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1622_inst_ack_0, ack => convTransposeA_CP_4108_elements(50)); -- 
    cr_4497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(50), ack => RPIPE_Block0_start_1622_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	54 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1622_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_Sample/rr
      -- 
    ca_4498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1622_inst_ack_1, ack => convTransposeA_CP_4108_elements(51)); -- 
    rr_4506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(51), ack => type_cast_1626_inst_req_0); -- 
    rr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(51), ack => RPIPE_Block0_start_1635_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_Sample/ra
      -- 
    ra_4507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_0, ack => convTransposeA_CP_4108_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	102 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1626_Update/$exit
      -- 
    ca_4512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_1, ack => convTransposeA_CP_4108_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_Update/cr
      -- CP-element group 54: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_sample_completed_
      -- 
    ra_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1635_inst_ack_0, ack => convTransposeA_CP_4108_elements(54)); -- 
    cr_4525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(54), ack => RPIPE_Block0_start_1635_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1635_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_Sample/rr
      -- 
    ca_4526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1635_inst_ack_1, ack => convTransposeA_CP_4108_elements(55)); -- 
    rr_4534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(55), ack => type_cast_1639_inst_req_0); -- 
    rr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(55), ack => RPIPE_Block0_start_1647_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_sample_completed_
      -- 
    ra_4535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1639_inst_ack_0, ack => convTransposeA_CP_4108_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	102 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1639_update_completed_
      -- 
    ca_4540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1639_inst_ack_1, ack => convTransposeA_CP_4108_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_Sample/ra
      -- 
    ra_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1647_inst_ack_0, ack => convTransposeA_CP_4108_elements(58)); -- 
    cr_4553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(58), ack => RPIPE_Block0_start_1647_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	62 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1647_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_Sample/rr
      -- 
    ca_4554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1647_inst_ack_1, ack => convTransposeA_CP_4108_elements(59)); -- 
    rr_4562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(59), ack => type_cast_1651_inst_req_0); -- 
    rr_4576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(59), ack => RPIPE_Block0_start_1660_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_Sample/ra
      -- CP-element group 60: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_Sample/$exit
      -- 
    ra_4563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1651_inst_ack_0, ack => convTransposeA_CP_4108_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	102 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1651_update_completed_
      -- 
    ca_4568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1651_inst_ack_1, ack => convTransposeA_CP_4108_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_sample_completed_
      -- 
    ra_4577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1660_inst_ack_0, ack => convTransposeA_CP_4108_elements(62)); -- 
    cr_4581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(62), ack => RPIPE_Block0_start_1660_inst_req_1); -- 
    -- CP-element group 63:  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1660_update_completed_
      -- 
    ca_4582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1660_inst_ack_1, ack => convTransposeA_CP_4108_elements(63)); -- 
    rr_4604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(63), ack => RPIPE_Block0_start_1672_inst_req_0); -- 
    rr_4590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(63), ack => type_cast_1664_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_Sample/ra
      -- CP-element group 64: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_sample_completed_
      -- 
    ra_4591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1664_inst_ack_0, ack => convTransposeA_CP_4108_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	102 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_Update/ca
      -- CP-element group 65: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1664_Update/$exit
      -- 
    ca_4596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1664_inst_ack_1, ack => convTransposeA_CP_4108_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_Sample/ra
      -- 
    ra_4605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1672_inst_ack_0, ack => convTransposeA_CP_4108_elements(66)); -- 
    cr_4609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(66), ack => RPIPE_Block0_start_1672_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1672_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_Sample/rr
      -- 
    ca_4610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1672_inst_ack_1, ack => convTransposeA_CP_4108_elements(67)); -- 
    rr_4618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(67), ack => type_cast_1676_inst_req_0); -- 
    rr_4632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(67), ack => RPIPE_Block0_start_1685_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_Sample/ra
      -- 
    ra_4619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1676_inst_ack_0, ack => convTransposeA_CP_4108_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	102 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1676_Update/ca
      -- 
    ca_4624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1676_inst_ack_1, ack => convTransposeA_CP_4108_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_update_start_
      -- 
    ra_4633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1685_inst_ack_0, ack => convTransposeA_CP_4108_elements(70)); -- 
    cr_4637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(70), ack => RPIPE_Block0_start_1685_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	74 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1685_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_Sample/rr
      -- 
    ca_4638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1685_inst_ack_1, ack => convTransposeA_CP_4108_elements(71)); -- 
    rr_4660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(71), ack => RPIPE_Block0_start_1703_inst_req_0); -- 
    rr_4646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(71), ack => type_cast_1689_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_sample_completed_
      -- 
    ra_4647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1689_inst_ack_0, ack => convTransposeA_CP_4108_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	102 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1689_Update/ca
      -- 
    ca_4652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1689_inst_ack_1, ack => convTransposeA_CP_4108_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	71 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_Update/cr
      -- 
    ra_4661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1703_inst_ack_0, ack => convTransposeA_CP_4108_elements(74)); -- 
    cr_4665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(74), ack => RPIPE_Block0_start_1703_inst_req_1); -- 
    -- CP-element group 75:  fork  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (9) 
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1703_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_Sample/rr
      -- 
    ca_4666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1703_inst_ack_1, ack => convTransposeA_CP_4108_elements(75)); -- 
    rr_4674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(75), ack => type_cast_1707_inst_req_0); -- 
    rr_4688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(75), ack => RPIPE_Block0_start_1721_inst_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_Sample/ra
      -- 
    ra_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1707_inst_ack_0, ack => convTransposeA_CP_4108_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	102 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1707_Update/ca
      -- 
    ca_4680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1707_inst_ack_1, ack => convTransposeA_CP_4108_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_update_start_
      -- CP-element group 78: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_Update/cr
      -- 
    ra_4689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1721_inst_ack_0, ack => convTransposeA_CP_4108_elements(78)); -- 
    cr_4693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(78), ack => RPIPE_Block0_start_1721_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1721_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_Sample/rr
      -- 
    ca_4694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1721_inst_ack_1, ack => convTransposeA_CP_4108_elements(79)); -- 
    rr_4716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(79), ack => RPIPE_Block0_start_1733_inst_req_0); -- 
    rr_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(79), ack => type_cast_1725_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_Sample/ra
      -- 
    ra_4703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1725_inst_ack_0, ack => convTransposeA_CP_4108_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	102 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1725_Update/ca
      -- 
    ca_4708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1725_inst_ack_1, ack => convTransposeA_CP_4108_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_Update/cr
      -- 
    ra_4717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1733_inst_ack_0, ack => convTransposeA_CP_4108_elements(82)); -- 
    cr_4721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(82), ack => RPIPE_Block0_start_1733_inst_req_1); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1733_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_Sample/rr
      -- 
    ca_4722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1733_inst_ack_1, ack => convTransposeA_CP_4108_elements(83)); -- 
    rr_4730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(83), ack => RPIPE_Block0_start_1736_inst_req_0); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_update_start_
      -- CP-element group 84: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_Update/cr
      -- 
    ra_4731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1736_inst_ack_0, ack => convTransposeA_CP_4108_elements(84)); -- 
    cr_4735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(84), ack => RPIPE_Block0_start_1736_inst_req_1); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1736_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_Sample/rr
      -- 
    ca_4736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1736_inst_ack_1, ack => convTransposeA_CP_4108_elements(85)); -- 
    rr_4744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(85), ack => RPIPE_Block0_start_1739_inst_req_0); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_update_start_
      -- CP-element group 86: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_Update/cr
      -- 
    ra_4745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1739_inst_ack_0, ack => convTransposeA_CP_4108_elements(86)); -- 
    cr_4749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(86), ack => RPIPE_Block0_start_1739_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	90 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1739_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_Sample/rr
      -- 
    ca_4750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1739_inst_ack_1, ack => convTransposeA_CP_4108_elements(87)); -- 
    rr_4758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(87), ack => type_cast_1743_inst_req_0); -- 
    rr_4772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(87), ack => RPIPE_Block0_start_1752_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_Sample/ra
      -- 
    ra_4759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1743_inst_ack_0, ack => convTransposeA_CP_4108_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	102 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1743_Update/ca
      -- 
    ca_4764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1743_inst_ack_1, ack => convTransposeA_CP_4108_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_update_start_
      -- CP-element group 90: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_Update/cr
      -- 
    ra_4773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1752_inst_ack_0, ack => convTransposeA_CP_4108_elements(90)); -- 
    cr_4777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(90), ack => RPIPE_Block0_start_1752_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1752_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_Sample/rr
      -- 
    ca_4778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1752_inst_ack_1, ack => convTransposeA_CP_4108_elements(91)); -- 
    rr_4786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(91), ack => type_cast_1756_inst_req_0); -- 
    rr_4800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(91), ack => RPIPE_Block0_start_1764_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_Sample/ra
      -- 
    ra_4787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1756_inst_ack_0, ack => convTransposeA_CP_4108_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	102 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1756_Update/ca
      -- 
    ca_4792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1756_inst_ack_1, ack => convTransposeA_CP_4108_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_Update/cr
      -- 
    ra_4801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1764_inst_ack_0, ack => convTransposeA_CP_4108_elements(94)); -- 
    cr_4805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(94), ack => RPIPE_Block0_start_1764_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1764_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_Sample/rr
      -- 
    ca_4806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1764_inst_ack_1, ack => convTransposeA_CP_4108_elements(95)); -- 
    rr_4814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(95), ack => type_cast_1768_inst_req_0); -- 
    rr_4828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(95), ack => RPIPE_Block0_start_1777_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_Sample/ra
      -- 
    ra_4815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_0, ack => convTransposeA_CP_4108_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	102 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1768_Update/ca
      -- 
    ca_4820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_1, ack => convTransposeA_CP_4108_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_Update/cr
      -- 
    ra_4829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1777_inst_ack_0, ack => convTransposeA_CP_4108_elements(98)); -- 
    cr_4833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(98), ack => RPIPE_Block0_start_1777_inst_req_1); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/RPIPE_Block0_start_1777_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_Sample/rr
      -- 
    ca_4834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1777_inst_ack_1, ack => convTransposeA_CP_4108_elements(99)); -- 
    rr_4842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(99), ack => type_cast_1781_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_Sample/ra
      -- 
    ra_4843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1781_inst_ack_0, ack => convTransposeA_CP_4108_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/type_cast_1781_Update/ca
      -- 
    ca_4848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1781_inst_ack_1, ack => convTransposeA_CP_4108_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	5 
    -- CP-element group 102: 	9 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	61 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	69 
    -- CP-element group 102: 	73 
    -- CP-element group 102: 	93 
    -- CP-element group 102: 	101 
    -- CP-element group 102: 	97 
    -- CP-element group 102: 	89 
    -- CP-element group 102: 	77 
    -- CP-element group 102: 	81 
    -- CP-element group 102: 	13 
    -- CP-element group 102: 	17 
    -- CP-element group 102: 	21 
    -- CP-element group 102: 	25 
    -- CP-element group 102: 	33 
    -- CP-element group 102: 	37 
    -- CP-element group 102: 	41 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	140 
    -- CP-element group 102: 	141 
    -- CP-element group 102: 	142 
    -- CP-element group 102: 	143 
    -- CP-element group 102:  members (16) 
      -- CP-element group 102: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787__exit__
      -- CP-element group 102: 	 branch_block_stmt_1482/assign_stmt_1794_to_assign_stmt_1816__entry__
      -- CP-element group 102: 	 branch_block_stmt_1482/assign_stmt_1794_to_assign_stmt_1816__exit__
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody
      -- CP-element group 102: 	 branch_block_stmt_1482/assign_stmt_1485_to_assign_stmt_1787/$exit
      -- CP-element group 102: 	 branch_block_stmt_1482/assign_stmt_1794_to_assign_stmt_1816/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/assign_stmt_1794_to_assign_stmt_1816/$exit
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1819/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1826/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1833/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1840/$entry
      -- CP-element group 102: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/$entry
      -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(5) & convTransposeA_CP_4108_elements(9) & convTransposeA_CP_4108_elements(57) & convTransposeA_CP_4108_elements(61) & convTransposeA_CP_4108_elements(53) & convTransposeA_CP_4108_elements(45) & convTransposeA_CP_4108_elements(65) & convTransposeA_CP_4108_elements(69) & convTransposeA_CP_4108_elements(73) & convTransposeA_CP_4108_elements(93) & convTransposeA_CP_4108_elements(101) & convTransposeA_CP_4108_elements(97) & convTransposeA_CP_4108_elements(89) & convTransposeA_CP_4108_elements(77) & convTransposeA_CP_4108_elements(81) & convTransposeA_CP_4108_elements(13) & convTransposeA_CP_4108_elements(17) & convTransposeA_CP_4108_elements(21) & convTransposeA_CP_4108_elements(25) & convTransposeA_CP_4108_elements(33) & convTransposeA_CP_4108_elements(37) & convTransposeA_CP_4108_elements(41);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	163 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_Sample/ra
      -- 
    ra_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_0, ack => convTransposeA_CP_4108_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	163 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	117 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_Update/ca
      -- 
    ca_4868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1881_inst_ack_1, ack => convTransposeA_CP_4108_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	163 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_Sample/ra
      -- 
    ra_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1885_inst_ack_0, ack => convTransposeA_CP_4108_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	163 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	117 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_Update/ca
      -- 
    ca_4882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1885_inst_ack_1, ack => convTransposeA_CP_4108_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	163 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_Sample/ra
      -- 
    ra_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1889_inst_ack_0, ack => convTransposeA_CP_4108_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	163 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	117 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_Update/ca
      -- 
    ca_4896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1889_inst_ack_1, ack => convTransposeA_CP_4108_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	163 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_Sample/ra
      -- 
    ra_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1919_inst_ack_0, ack => convTransposeA_CP_4108_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	163 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (16) 
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_resized_1
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_scaled_1
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_computed_1
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_resize_1/$entry
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_resize_1/$exit
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_resize_1/index_resize_req
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_resize_1/index_resize_ack
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_scale_1/$entry
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_scale_1/$exit
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_scale_1/scale_rename_req
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_index_scale_1/scale_rename_ack
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_Sample/req
      -- 
    ca_4910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1919_inst_ack_1, ack => convTransposeA_CP_4108_elements(110)); -- 
    req_4935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(110), ack => array_obj_ref_1925_index_offset_req_0); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	127 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_sample_complete
      -- CP-element group 111: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_Sample/ack
      -- 
    ack_4936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1925_index_offset_ack_0, ack => convTransposeA_CP_4108_elements(111)); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	163 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (11) 
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_root_address_calculated
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_offset_calculated
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_Update/ack
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_base_plus_offset/$entry
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_base_plus_offset/$exit
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_base_plus_offset/sum_rename_req
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_base_plus_offset/sum_rename_ack
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_request/$entry
      -- CP-element group 112: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_request/req
      -- 
    ack_4941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1925_index_offset_ack_1, ack => convTransposeA_CP_4108_elements(112)); -- 
    req_4950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(112), ack => addr_of_1926_final_reg_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_request/$exit
      -- CP-element group 113: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_request/ack
      -- 
    ack_4951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1926_final_reg_ack_0, ack => convTransposeA_CP_4108_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	163 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (24) 
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_complete/$exit
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_complete/ack
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_address_calculated
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_word_address_calculated
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_root_address_calculated
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_address_resized
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_addr_resize/$entry
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_addr_resize/$exit
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_addr_resize/base_resize_req
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_addr_resize/base_resize_ack
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_plus_offset/$entry
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_plus_offset/$exit
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_plus_offset/sum_rename_req
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_base_plus_offset/sum_rename_ack
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_word_addrgen/$entry
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_word_addrgen/$exit
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_word_addrgen/root_register_req
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_word_addrgen/root_register_ack
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Sample/word_access_start/$entry
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Sample/word_access_start/word_0/$entry
      -- CP-element group 114: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Sample/word_access_start/word_0/rr
      -- 
    ack_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1926_final_reg_ack_1, ack => convTransposeA_CP_4108_elements(114)); -- 
    rr_4989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(114), ack => ptr_deref_1930_load_0_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Sample/word_access_start/$exit
      -- CP-element group 115: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Sample/word_access_start/word_0/$exit
      -- CP-element group 115: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Sample/word_access_start/word_0/ra
      -- 
    ra_4990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1930_load_0_ack_0, ack => convTransposeA_CP_4108_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	163 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	122 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/word_access_complete/$exit
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/word_access_complete/word_0/$exit
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/word_access_complete/word_0/ca
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/ptr_deref_1930_Merge/$entry
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/ptr_deref_1930_Merge/$exit
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/ptr_deref_1930_Merge/merge_req
      -- CP-element group 116: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/ptr_deref_1930_Merge/merge_ack
      -- 
    ca_5001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1930_load_0_ack_1, ack => convTransposeA_CP_4108_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	108 
    -- CP-element group 117: 	104 
    -- CP-element group 117: 	106 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (13) 
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_resized_1
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_scaled_1
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_computed_1
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_resize_1/$entry
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_resize_1/$exit
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_resize_1/index_resize_req
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_resize_1/index_resize_ack
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_scale_1/$entry
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_scale_1/$exit
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_scale_1/scale_rename_req
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_index_scale_1/scale_rename_ack
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_Sample/req
      -- 
    req_5031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(117), ack => array_obj_ref_1948_index_offset_req_0); -- 
    convTransposeA_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(108) & convTransposeA_CP_4108_elements(104) & convTransposeA_CP_4108_elements(106);
      gj_convTransposeA_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	127 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_sample_complete
      -- CP-element group 118: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_Sample/ack
      -- 
    ack_5032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1948_index_offset_ack_0, ack => convTransposeA_CP_4108_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	163 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (11) 
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_offset_calculated
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_Update/ack
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_request/$entry
      -- CP-element group 119: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_request/req
      -- 
    ack_5037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1948_index_offset_ack_1, ack => convTransposeA_CP_4108_elements(119)); -- 
    req_5046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(119), ack => addr_of_1949_final_reg_req_0); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_request/$exit
      -- CP-element group 120: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_request/ack
      -- 
    ack_5047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1949_final_reg_ack_0, ack => convTransposeA_CP_4108_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	163 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (19) 
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_complete/$exit
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_complete/ack
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_word_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_root_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_address_resized
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_addr_resize/$entry
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_addr_resize/$exit
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_addr_resize/base_resize_req
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_addr_resize/base_resize_ack
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_plus_offset/$entry
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_plus_offset/$exit
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_plus_offset/sum_rename_req
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_base_plus_offset/sum_rename_ack
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_word_addrgen/$entry
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_word_addrgen/$exit
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_word_addrgen/root_register_req
      -- CP-element group 121: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_word_addrgen/root_register_ack
      -- 
    ack_5052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1949_final_reg_ack_1, ack => convTransposeA_CP_4108_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: 	116 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (9) 
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/ptr_deref_1952_Split/$entry
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/ptr_deref_1952_Split/$exit
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/ptr_deref_1952_Split/split_req
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/ptr_deref_1952_Split/split_ack
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/word_access_start/$entry
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/word_access_start/word_0/$entry
      -- CP-element group 122: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/word_access_start/word_0/rr
      -- 
    rr_5090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(122), ack => ptr_deref_1952_store_0_req_0); -- 
    convTransposeA_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(121) & convTransposeA_CP_4108_elements(116);
      gj_convTransposeA_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (5) 
      -- CP-element group 123: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/word_access_start/$exit
      -- CP-element group 123: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/word_access_start/word_0/$exit
      -- CP-element group 123: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Sample/word_access_start/word_0/ra
      -- 
    ra_5091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1952_store_0_ack_0, ack => convTransposeA_CP_4108_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	163 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Update/word_access_complete/$exit
      -- CP-element group 124: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Update/word_access_complete/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Update/word_access_complete/word_0/ca
      -- 
    ca_5102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1952_store_0_ack_1, ack => convTransposeA_CP_4108_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	163 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_Sample/ra
      -- 
    ra_5111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_0, ack => convTransposeA_CP_4108_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	163 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_Update/ca
      -- 
    ca_5116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_1, ack => convTransposeA_CP_4108_elements(126)); -- 
    -- CP-element group 127:  branch  join  transition  place  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	118 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	126 
    -- CP-element group 127: 	111 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (10) 
      -- CP-element group 127: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969__exit__
      -- CP-element group 127: 	 branch_block_stmt_1482/if_stmt_1970__entry__
      -- CP-element group 127: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/$exit
      -- CP-element group 127: 	 branch_block_stmt_1482/if_stmt_1970_dead_link/$entry
      -- CP-element group 127: 	 branch_block_stmt_1482/if_stmt_1970_eval_test/$entry
      -- CP-element group 127: 	 branch_block_stmt_1482/if_stmt_1970_eval_test/$exit
      -- CP-element group 127: 	 branch_block_stmt_1482/if_stmt_1970_eval_test/branch_req
      -- CP-element group 127: 	 branch_block_stmt_1482/R_cmp_1971_place
      -- CP-element group 127: 	 branch_block_stmt_1482/if_stmt_1970_if_link/$entry
      -- CP-element group 127: 	 branch_block_stmt_1482/if_stmt_1970_else_link/$entry
      -- 
    branch_req_5124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(127), ack => if_stmt_1970_branch_req_0); -- 
    convTransposeA_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(118) & convTransposeA_CP_4108_elements(124) & convTransposeA_CP_4108_elements(126) & convTransposeA_CP_4108_elements(111);
      gj_convTransposeA_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	178 
    -- CP-element group 128: 	179 
    -- CP-element group 128: 	172 
    -- CP-element group 128: 	173 
    -- CP-element group 128: 	175 
    -- CP-element group 128: 	176 
    -- CP-element group 128:  members (40) 
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/merge_stmt_1976__exit__
      -- CP-element group 128: 	 branch_block_stmt_1482/assign_stmt_1982__entry__
      -- CP-element group 128: 	 branch_block_stmt_1482/assign_stmt_1982__exit__
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_1482/if_stmt_1970_if_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_1482/if_stmt_1970_if_link/if_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/whilex_xbody_ifx_xthen
      -- CP-element group 128: 	 branch_block_stmt_1482/assign_stmt_1982/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/assign_stmt_1982/$exit
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 128: 	 branch_block_stmt_1482/merge_stmt_1976_PhiReqMerge
      -- CP-element group 128: 	 branch_block_stmt_1482/merge_stmt_1976_PhiAck/$entry
      -- CP-element group 128: 	 branch_block_stmt_1482/merge_stmt_1976_PhiAck/$exit
      -- CP-element group 128: 	 branch_block_stmt_1482/merge_stmt_1976_PhiAck/dummy
      -- 
    if_choice_transition_5129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1970_branch_ack_1, ack => convTransposeA_CP_4108_elements(128)); -- 
    cr_5465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(128), ack => type_cast_2050_inst_req_1); -- 
    rr_5460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(128), ack => type_cast_2050_inst_req_0); -- 
    cr_5511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(128), ack => type_cast_2035_inst_req_1); -- 
    cr_5488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(128), ack => type_cast_2042_inst_req_1); -- 
    rr_5483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(128), ack => type_cast_2042_inst_req_0); -- 
    rr_5506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(128), ack => type_cast_2035_inst_req_0); -- 
    -- CP-element group 129:  fork  transition  place  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: 	131 
    -- CP-element group 129: 	133 
    -- CP-element group 129: 	135 
    -- CP-element group 129:  members (24) 
      -- CP-element group 129: 	 branch_block_stmt_1482/merge_stmt_1984__exit__
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024__entry__
      -- CP-element group 129: 	 branch_block_stmt_1482/if_stmt_1970_else_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_1482/if_stmt_1970_else_link/else_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_1482/whilex_xbody_ifx_xelse
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/$entry
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_update_start_
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_Sample/rr
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_update_start_
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_update_start_
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_1482/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_1482/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 129: 	 branch_block_stmt_1482/merge_stmt_1984_PhiReqMerge
      -- CP-element group 129: 	 branch_block_stmt_1482/merge_stmt_1984_PhiAck/$entry
      -- CP-element group 129: 	 branch_block_stmt_1482/merge_stmt_1984_PhiAck/$exit
      -- CP-element group 129: 	 branch_block_stmt_1482/merge_stmt_1984_PhiAck/dummy
      -- 
    else_choice_transition_5133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1970_branch_ack_0, ack => convTransposeA_CP_4108_elements(129)); -- 
    rr_5149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(129), ack => type_cast_1993_inst_req_0); -- 
    cr_5154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(129), ack => type_cast_1993_inst_req_1); -- 
    cr_5168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(129), ack => type_cast_2002_inst_req_1); -- 
    cr_5182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(129), ack => type_cast_2018_inst_req_1); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_Sample/ra
      -- 
    ra_5150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_0, ack => convTransposeA_CP_4108_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_1993_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_Sample/rr
      -- 
    ca_5155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_1, ack => convTransposeA_CP_4108_elements(131)); -- 
    rr_5163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(131), ack => type_cast_2002_inst_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_Sample/ra
      -- 
    ra_5164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2002_inst_ack_0, ack => convTransposeA_CP_4108_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	129 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2002_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_Sample/rr
      -- 
    ca_5169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2002_inst_ack_1, ack => convTransposeA_CP_4108_elements(133)); -- 
    rr_5177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(133), ack => type_cast_2018_inst_req_0); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_Sample/ra
      -- 
    ra_5178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2018_inst_ack_0, ack => convTransposeA_CP_4108_elements(134)); -- 
    -- CP-element group 135:  branch  transition  place  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	129 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (13) 
      -- CP-element group 135: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024__exit__
      -- CP-element group 135: 	 branch_block_stmt_1482/if_stmt_2025__entry__
      -- CP-element group 135: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/$exit
      -- CP-element group 135: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1482/assign_stmt_1990_to_assign_stmt_2024/type_cast_2018_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_1482/if_stmt_2025_dead_link/$entry
      -- CP-element group 135: 	 branch_block_stmt_1482/if_stmt_2025_eval_test/$entry
      -- CP-element group 135: 	 branch_block_stmt_1482/if_stmt_2025_eval_test/$exit
      -- CP-element group 135: 	 branch_block_stmt_1482/if_stmt_2025_eval_test/branch_req
      -- CP-element group 135: 	 branch_block_stmt_1482/R_cmp238_2026_place
      -- CP-element group 135: 	 branch_block_stmt_1482/if_stmt_2025_if_link/$entry
      -- CP-element group 135: 	 branch_block_stmt_1482/if_stmt_2025_else_link/$entry
      -- 
    ca_5183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2018_inst_ack_1, ack => convTransposeA_CP_4108_elements(135)); -- 
    branch_req_5191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(135), ack => if_stmt_2025_branch_req_0); -- 
    -- CP-element group 136:  transition  place  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (15) 
      -- CP-element group 136: 	 branch_block_stmt_1482/merge_stmt_2059__exit__
      -- CP-element group 136: 	 branch_block_stmt_1482/assign_stmt_2064__entry__
      -- CP-element group 136: 	 branch_block_stmt_1482/merge_stmt_2059_PhiAck/dummy
      -- CP-element group 136: 	 branch_block_stmt_1482/merge_stmt_2059_PhiAck/$exit
      -- CP-element group 136: 	 branch_block_stmt_1482/merge_stmt_2059_PhiAck/$entry
      -- CP-element group 136: 	 branch_block_stmt_1482/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 136: 	 branch_block_stmt_1482/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 136: 	 branch_block_stmt_1482/merge_stmt_2059_PhiReqMerge
      -- CP-element group 136: 	 branch_block_stmt_1482/if_stmt_2025_if_link/$exit
      -- CP-element group 136: 	 branch_block_stmt_1482/if_stmt_2025_if_link/if_choice_transition
      -- CP-element group 136: 	 branch_block_stmt_1482/ifx_xelse_whilex_xend
      -- CP-element group 136: 	 branch_block_stmt_1482/assign_stmt_2064/$entry
      -- CP-element group 136: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_Sample/req
      -- 
    if_choice_transition_5196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2025_branch_ack_1, ack => convTransposeA_CP_4108_elements(136)); -- 
    req_5216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(136), ack => WPIPE_Block0_done_2061_inst_req_0); -- 
    -- CP-element group 137:  fork  transition  place  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	164 
    -- CP-element group 137: 	165 
    -- CP-element group 137: 	167 
    -- CP-element group 137: 	168 
    -- CP-element group 137: 	170 
    -- CP-element group 137:  members (22) 
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/Sample/rr
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/Sample/rr
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/Update/cr
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2032/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/Update/cr
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1482/if_stmt_2025_else_link/$exit
      -- CP-element group 137: 	 branch_block_stmt_1482/if_stmt_2025_else_link/else_choice_transition
      -- CP-element group 137: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249
      -- 
    else_choice_transition_5200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2025_branch_ack_0, ack => convTransposeA_CP_4108_elements(137)); -- 
    rr_5426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(137), ack => type_cast_2044_inst_req_0); -- 
    rr_5403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(137), ack => type_cast_2048_inst_req_0); -- 
    cr_5408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(137), ack => type_cast_2048_inst_req_1); -- 
    cr_5431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(137), ack => type_cast_2044_inst_req_1); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_update_start_
      -- CP-element group 138: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_Sample/ack
      -- CP-element group 138: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_Update/req
      -- 
    ack_5217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_2061_inst_ack_0, ack => convTransposeA_CP_4108_elements(138)); -- 
    req_5221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(138), ack => WPIPE_Block0_done_2061_inst_req_1); -- 
    -- CP-element group 139:  transition  place  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (16) 
      -- CP-element group 139: 	 $exit
      -- CP-element group 139: 	 branch_block_stmt_1482/$exit
      -- CP-element group 139: 	 branch_block_stmt_1482/branch_block_stmt_1482__exit__
      -- CP-element group 139: 	 branch_block_stmt_1482/assign_stmt_2064__exit__
      -- CP-element group 139: 	 branch_block_stmt_1482/return__
      -- CP-element group 139: 	 branch_block_stmt_1482/merge_stmt_2066__exit__
      -- CP-element group 139: 	 branch_block_stmt_1482/merge_stmt_2066_PhiReqMerge
      -- CP-element group 139: 	 branch_block_stmt_1482/merge_stmt_2066_PhiAck/dummy
      -- CP-element group 139: 	 branch_block_stmt_1482/merge_stmt_2066_PhiAck/$exit
      -- CP-element group 139: 	 branch_block_stmt_1482/merge_stmt_2066_PhiAck/$entry
      -- CP-element group 139: 	 branch_block_stmt_1482/return___PhiReq/$exit
      -- CP-element group 139: 	 branch_block_stmt_1482/return___PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_1482/assign_stmt_2064/$exit
      -- CP-element group 139: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_1482/assign_stmt_2064/WPIPE_Block0_done_2061_Update/ack
      -- 
    ack_5222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_2061_inst_ack_1, ack => convTransposeA_CP_4108_elements(139)); -- 
    -- CP-element group 140:  transition  output  delay-element  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	102 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	144 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1819/$exit
      -- CP-element group 140: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/$exit
      -- CP-element group 140: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1823_konst_delay_trans
      -- CP-element group 140: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_req
      -- 
    phi_stmt_1819_req_5233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1819_req_5233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(140), ack => phi_stmt_1819_req_0); -- 
    -- Element group convTransposeA_CP_4108_elements(140) is a control-delay.
    cp_element_140_delay: control_delay_element  generic map(name => " 140_delay", delay_value => 1)  port map(req => convTransposeA_CP_4108_elements(102), ack => convTransposeA_CP_4108_elements(140), clk => clk, reset =>reset);
    -- CP-element group 141:  transition  output  delay-element  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	102 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	144 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1826/$exit
      -- CP-element group 141: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/$exit
      -- CP-element group 141: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1830_konst_delay_trans
      -- CP-element group 141: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_req
      -- 
    phi_stmt_1826_req_5241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1826_req_5241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(141), ack => phi_stmt_1826_req_0); -- 
    -- Element group convTransposeA_CP_4108_elements(141) is a control-delay.
    cp_element_141_delay: control_delay_element  generic map(name => " 141_delay", delay_value => 1)  port map(req => convTransposeA_CP_4108_elements(102), ack => convTransposeA_CP_4108_elements(141), clk => clk, reset =>reset);
    -- CP-element group 142:  transition  output  delay-element  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	102 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1833/$exit
      -- CP-element group 142: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/$exit
      -- CP-element group 142: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1837_konst_delay_trans
      -- CP-element group 142: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_req
      -- 
    phi_stmt_1833_req_5249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1833_req_5249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(142), ack => phi_stmt_1833_req_0); -- 
    -- Element group convTransposeA_CP_4108_elements(142) is a control-delay.
    cp_element_142_delay: control_delay_element  generic map(name => " 142_delay", delay_value => 1)  port map(req => convTransposeA_CP_4108_elements(102), ack => convTransposeA_CP_4108_elements(142), clk => clk, reset =>reset);
    -- CP-element group 143:  transition  output  delay-element  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	102 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1840/$exit
      -- CP-element group 143: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/$exit
      -- CP-element group 143: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1844_konst_delay_trans
      -- CP-element group 143: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_req
      -- 
    phi_stmt_1840_req_5257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1840_req_5257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(143), ack => phi_stmt_1840_req_0); -- 
    -- Element group convTransposeA_CP_4108_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => convTransposeA_CP_4108_elements(102), ack => convTransposeA_CP_4108_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  join  transition  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	140 
    -- CP-element group 144: 	141 
    -- CP-element group 144: 	142 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	158 
    -- CP-element group 144:  members (1) 
      -- CP-element group 144: 	 branch_block_stmt_1482/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(140) & convTransposeA_CP_4108_elements(141) & convTransposeA_CP_4108_elements(142) & convTransposeA_CP_4108_elements(143);
      gj_convTransposeA_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	1 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/Sample/ra
      -- 
    ra_5277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_0, ack => convTransposeA_CP_4108_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	1 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/Update/ca
      -- 
    ca_5282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_1, ack => convTransposeA_CP_4108_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	157 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/$exit
      -- CP-element group 147: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/$exit
      -- CP-element group 147: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/$exit
      -- CP-element group 147: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_sources/type_cast_1825/SplitProtocol/$exit
      -- CP-element group 147: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1819/phi_stmt_1819_req
      -- 
    phi_stmt_1819_req_5283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1819_req_5283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(147), ack => phi_stmt_1819_req_1); -- 
    convTransposeA_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(145) & convTransposeA_CP_4108_elements(146);
      gj_convTransposeA_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	1 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/Sample/ra
      -- 
    ra_5300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_0, ack => convTransposeA_CP_4108_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	1 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/Update/ca
      -- 
    ca_5305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1832_inst_ack_1, ack => convTransposeA_CP_4108_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	157 
    -- CP-element group 150:  members (5) 
      -- CP-element group 150: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/$exit
      -- CP-element group 150: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/$exit
      -- CP-element group 150: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/$exit
      -- CP-element group 150: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_sources/type_cast_1832/SplitProtocol/$exit
      -- CP-element group 150: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1826/phi_stmt_1826_req
      -- 
    phi_stmt_1826_req_5306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1826_req_5306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(150), ack => phi_stmt_1826_req_1); -- 
    convTransposeA_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(148) & convTransposeA_CP_4108_elements(149);
      gj_convTransposeA_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	1 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (2) 
      -- CP-element group 151: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/Sample/ra
      -- 
    ra_5323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1839_inst_ack_0, ack => convTransposeA_CP_4108_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	1 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/Update/ca
      -- 
    ca_5328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1839_inst_ack_1, ack => convTransposeA_CP_4108_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	157 
    -- CP-element group 153:  members (5) 
      -- CP-element group 153: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/$exit
      -- CP-element group 153: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/$exit
      -- CP-element group 153: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/$exit
      -- CP-element group 153: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_sources/type_cast_1839/SplitProtocol/$exit
      -- CP-element group 153: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1833/phi_stmt_1833_req
      -- 
    phi_stmt_1833_req_5329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1833_req_5329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(153), ack => phi_stmt_1833_req_1); -- 
    convTransposeA_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(151) & convTransposeA_CP_4108_elements(152);
      gj_convTransposeA_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	1 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (2) 
      -- CP-element group 154: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/Sample/ra
      -- 
    ra_5346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1846_inst_ack_0, ack => convTransposeA_CP_4108_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	1 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (2) 
      -- CP-element group 155: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/Update/ca
      -- 
    ca_5351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1846_inst_ack_1, ack => convTransposeA_CP_4108_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/$exit
      -- CP-element group 156: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/$exit
      -- CP-element group 156: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/$exit
      -- CP-element group 156: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_sources/type_cast_1846/SplitProtocol/$exit
      -- CP-element group 156: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/phi_stmt_1840/phi_stmt_1840_req
      -- 
    phi_stmt_1840_req_5352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1840_req_5352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(156), ack => phi_stmt_1840_req_1); -- 
    convTransposeA_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(154) & convTransposeA_CP_4108_elements(155);
      gj_convTransposeA_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	147 
    -- CP-element group 157: 	150 
    -- CP-element group 157: 	153 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1482/ifx_xend249_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(147) & convTransposeA_CP_4108_elements(150) & convTransposeA_CP_4108_elements(153) & convTransposeA_CP_4108_elements(156);
      gj_convTransposeA_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  merge  fork  transition  place  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	144 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	160 
    -- CP-element group 158: 	161 
    -- CP-element group 158: 	162 
    -- CP-element group 158:  members (2) 
      -- CP-element group 158: 	 branch_block_stmt_1482/merge_stmt_1818_PhiReqMerge
      -- CP-element group 158: 	 branch_block_stmt_1482/merge_stmt_1818_PhiAck/$entry
      -- 
    convTransposeA_CP_4108_elements(158) <= OrReduce(convTransposeA_CP_4108_elements(144) & convTransposeA_CP_4108_elements(157));
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	163 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1482/merge_stmt_1818_PhiAck/phi_stmt_1819_ack
      -- 
    phi_stmt_1819_ack_5357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1819_ack_0, ack => convTransposeA_CP_4108_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	163 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_1482/merge_stmt_1818_PhiAck/phi_stmt_1826_ack
      -- 
    phi_stmt_1826_ack_5358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1826_ack_0, ack => convTransposeA_CP_4108_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	158 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1482/merge_stmt_1818_PhiAck/phi_stmt_1833_ack
      -- 
    phi_stmt_1833_ack_5359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1833_ack_0, ack => convTransposeA_CP_4108_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	158 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_1482/merge_stmt_1818_PhiAck/phi_stmt_1840_ack
      -- 
    phi_stmt_1840_ack_5360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1840_ack_0, ack => convTransposeA_CP_4108_elements(162)); -- 
    -- CP-element group 163:  join  fork  transition  place  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	159 
    -- CP-element group 163: 	160 
    -- CP-element group 163: 	161 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	119 
    -- CP-element group 163: 	121 
    -- CP-element group 163: 	124 
    -- CP-element group 163: 	125 
    -- CP-element group 163: 	126 
    -- CP-element group 163: 	112 
    -- CP-element group 163: 	116 
    -- CP-element group 163: 	114 
    -- CP-element group 163: 	108 
    -- CP-element group 163: 	109 
    -- CP-element group 163: 	110 
    -- CP-element group 163: 	103 
    -- CP-element group 163: 	104 
    -- CP-element group 163: 	105 
    -- CP-element group 163: 	106 
    -- CP-element group 163: 	107 
    -- CP-element group 163:  members (56) 
      -- CP-element group 163: 	 branch_block_stmt_1482/merge_stmt_1818__exit__
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969__entry__
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1881_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1885_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1889_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1919_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_update_start
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1925_final_index_sum_regn_Update/req
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1926_complete/req
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/word_access_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/word_access_complete/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1930_Update/word_access_complete/word_0/cr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_update_start
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/array_obj_ref_1948_final_index_sum_regn_Update/req
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/addr_of_1949_complete/req
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Update/word_access_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Update/word_access_complete/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/ptr_deref_1952_Update/word_access_complete/word_0/cr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1482/assign_stmt_1853_to_assign_stmt_1969/type_cast_1957_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_1482/merge_stmt_1818_PhiAck/$exit
      -- 
    rr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1881_inst_req_0); -- 
    cr_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1881_inst_req_1); -- 
    rr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1885_inst_req_0); -- 
    cr_4881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1885_inst_req_1); -- 
    rr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1889_inst_req_0); -- 
    cr_4895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1889_inst_req_1); -- 
    rr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1919_inst_req_0); -- 
    cr_4909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1919_inst_req_1); -- 
    req_4940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => array_obj_ref_1925_index_offset_req_1); -- 
    req_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => addr_of_1926_final_reg_req_1); -- 
    cr_5000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => ptr_deref_1930_load_0_req_1); -- 
    req_5036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => array_obj_ref_1948_index_offset_req_1); -- 
    req_5051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => addr_of_1949_final_reg_req_1); -- 
    cr_5101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => ptr_deref_1952_store_0_req_1); -- 
    rr_5110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1957_inst_req_0); -- 
    cr_5115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(163), ack => type_cast_1957_inst_req_1); -- 
    convTransposeA_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(159) & convTransposeA_CP_4108_elements(160) & convTransposeA_CP_4108_elements(161) & convTransposeA_CP_4108_elements(162);
      gj_convTransposeA_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	137 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/Sample/ra
      -- 
    ra_5404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2048_inst_ack_0, ack => convTransposeA_CP_4108_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	137 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/Update/ca
      -- CP-element group 165: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/Update/$exit
      -- 
    ca_5409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2048_inst_ack_1, ack => convTransposeA_CP_4108_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	171 
    -- CP-element group 166:  members (5) 
      -- CP-element group 166: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_req
      -- CP-element group 166: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/$exit
      -- CP-element group 166: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/SplitProtocol/$exit
      -- CP-element group 166: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2048/$exit
      -- CP-element group 166: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/$exit
      -- 
    phi_stmt_2045_req_5410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2045_req_5410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(166), ack => phi_stmt_2045_req_0); -- 
    convTransposeA_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(164) & convTransposeA_CP_4108_elements(165);
      gj_convTransposeA_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	137 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/Sample/$exit
      -- 
    ra_5427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2044_inst_ack_0, ack => convTransposeA_CP_4108_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	137 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (2) 
      -- CP-element group 168: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/Update/ca
      -- 
    ca_5432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2044_inst_ack_1, ack => convTransposeA_CP_4108_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (5) 
      -- CP-element group 169: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/$exit
      -- CP-element group 169: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/$exit
      -- CP-element group 169: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/SplitProtocol/$exit
      -- CP-element group 169: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_req
      -- CP-element group 169: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2044/$exit
      -- 
    phi_stmt_2039_req_5433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2039_req_5433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(169), ack => phi_stmt_2039_req_1); -- 
    convTransposeA_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(167) & convTransposeA_CP_4108_elements(168);
      gj_convTransposeA_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  transition  output  delay-element  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	137 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_req
      -- CP-element group 170: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2038_konst_delay_trans
      -- CP-element group 170: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/$exit
      -- CP-element group 170: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/phi_stmt_2032/$exit
      -- 
    phi_stmt_2032_req_5441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2032_req_5441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(170), ack => phi_stmt_2032_req_1); -- 
    -- Element group convTransposeA_CP_4108_elements(170) is a control-delay.
    cp_element_170_delay: control_delay_element  generic map(name => " 170_delay", delay_value => 1)  port map(req => convTransposeA_CP_4108_elements(137), ack => convTransposeA_CP_4108_elements(170), clk => clk, reset =>reset);
    -- CP-element group 171:  join  transition  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	166 
    -- CP-element group 171: 	169 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	182 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 branch_block_stmt_1482/ifx_xelse_ifx_xend249_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(166) & convTransposeA_CP_4108_elements(169) & convTransposeA_CP_4108_elements(170);
      gj_convTransposeA_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	128 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/Sample/ra
      -- CP-element group 172: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/Sample/$exit
      -- 
    ra_5461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2050_inst_ack_0, ack => convTransposeA_CP_4108_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	128 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (2) 
      -- CP-element group 173: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/Update/ca
      -- CP-element group 173: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/Update/$exit
      -- 
    ca_5466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2050_inst_ack_1, ack => convTransposeA_CP_4108_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	181 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_req
      -- CP-element group 174: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/SplitProtocol/$exit
      -- CP-element group 174: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/type_cast_2050/$exit
      -- CP-element group 174: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/phi_stmt_2045_sources/$exit
      -- CP-element group 174: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2045/$exit
      -- 
    phi_stmt_2045_req_5467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2045_req_5467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(174), ack => phi_stmt_2045_req_1); -- 
    convTransposeA_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(172) & convTransposeA_CP_4108_elements(173);
      gj_convTransposeA_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	128 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (2) 
      -- CP-element group 175: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/Sample/ra
      -- 
    ra_5484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2042_inst_ack_0, ack => convTransposeA_CP_4108_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	128 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/Update/ca
      -- CP-element group 176: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/Update/$exit
      -- 
    ca_5489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2042_inst_ack_1, ack => convTransposeA_CP_4108_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	181 
    -- CP-element group 177:  members (5) 
      -- CP-element group 177: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/$exit
      -- CP-element group 177: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/type_cast_2042/SplitProtocol/$exit
      -- CP-element group 177: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_sources/$exit
      -- CP-element group 177: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/$exit
      -- CP-element group 177: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2039/phi_stmt_2039_req
      -- 
    phi_stmt_2039_req_5490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2039_req_5490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(177), ack => phi_stmt_2039_req_0); -- 
    convTransposeA_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(175) & convTransposeA_CP_4108_elements(176);
      gj_convTransposeA_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	128 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/Sample/ra
      -- CP-element group 178: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/Sample/$exit
      -- 
    ra_5507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2035_inst_ack_0, ack => convTransposeA_CP_4108_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	128 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/Update/ca
      -- CP-element group 179: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/Update/$exit
      -- 
    ca_5512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2035_inst_ack_1, ack => convTransposeA_CP_4108_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (5) 
      -- CP-element group 180: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/$exit
      -- CP-element group 180: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/$exit
      -- CP-element group 180: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/$exit
      -- CP-element group 180: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_req
      -- CP-element group 180: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/phi_stmt_2032/phi_stmt_2032_sources/type_cast_2035/SplitProtocol/$exit
      -- 
    phi_stmt_2032_req_5513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2032_req_5513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4108_elements(180), ack => phi_stmt_2032_req_0); -- 
    convTransposeA_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(178) & convTransposeA_CP_4108_elements(179);
      gj_convTransposeA_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: 	174 
    -- CP-element group 181: 	177 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_1482/ifx_xthen_ifx_xend249_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(180) & convTransposeA_CP_4108_elements(174) & convTransposeA_CP_4108_elements(177);
      gj_convTransposeA_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  merge  fork  transition  place  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	171 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_1482/merge_stmt_2031_PhiAck/$entry
      -- CP-element group 182: 	 branch_block_stmt_1482/merge_stmt_2031_PhiReqMerge
      -- 
    convTransposeA_CP_4108_elements(182) <= OrReduce(convTransposeA_CP_4108_elements(171) & convTransposeA_CP_4108_elements(181));
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	186 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_1482/merge_stmt_2031_PhiAck/phi_stmt_2032_ack
      -- 
    phi_stmt_2032_ack_5518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2032_ack_0, ack => convTransposeA_CP_4108_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_1482/merge_stmt_2031_PhiAck/phi_stmt_2039_ack
      -- 
    phi_stmt_2039_ack_5519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2039_ack_0, ack => convTransposeA_CP_4108_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_1482/merge_stmt_2031_PhiAck/phi_stmt_2045_ack
      -- 
    phi_stmt_2045_ack_5520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2045_ack_0, ack => convTransposeA_CP_4108_elements(185)); -- 
    -- CP-element group 186:  join  transition  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	183 
    -- CP-element group 186: 	184 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	1 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_1482/merge_stmt_2031_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_4108_elements(183) & convTransposeA_CP_4108_elements(184) & convTransposeA_CP_4108_elements(185);
      gj_convTransposeA_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4108_elements(186), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom207_1947_resized : std_logic_vector(13 downto 0);
    signal R_idxprom207_1947_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1924_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1924_scaled : std_logic_vector(13 downto 0);
    signal add103_1695 : std_logic_vector(31 downto 0);
    signal add108_1713 : std_logic_vector(31 downto 0);
    signal add113_1731 : std_logic_vector(31 downto 0);
    signal add135_1762 : std_logic_vector(63 downto 0);
    signal add147_1787 : std_logic_vector(63 downto 0);
    signal add167_1794 : std_logic_vector(15 downto 0);
    signal add16_1532 : std_logic_vector(31 downto 0);
    signal add180_1805 : std_logic_vector(15 downto 0);
    signal add199_1900 : std_logic_vector(63 downto 0);
    signal add201_1910 : std_logic_vector(63 downto 0);
    signal add212_1964 : std_logic_vector(31 downto 0);
    signal add219_1982 : std_logic_vector(15 downto 0);
    signal add28_1557 : std_logic_vector(31 downto 0);
    signal add52_1589 : std_logic_vector(15 downto 0);
    signal add64_1614 : std_logic_vector(15 downto 0);
    signal add86_1645 : std_logic_vector(15 downto 0);
    signal add95_1670 : std_logic_vector(15 downto 0);
    signal add_1507 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1858 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1925_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1925_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1948_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1948_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1948_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1948_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1948_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1948_root_address : std_logic_vector(13 downto 0);
    signal arrayidx203_1927 : std_logic_vector(31 downto 0);
    signal arrayidx208_1950 : std_logic_vector(31 downto 0);
    signal call101_1686 : std_logic_vector(7 downto 0);
    signal call106_1704 : std_logic_vector(7 downto 0);
    signal call111_1722 : std_logic_vector(7 downto 0);
    signal call114_1734 : std_logic_vector(7 downto 0);
    signal call121_1737 : std_logic_vector(7 downto 0);
    signal call126_1740 : std_logic_vector(7 downto 0);
    signal call133_1753 : std_logic_vector(7 downto 0);
    signal call138_1765 : std_logic_vector(7 downto 0);
    signal call145_1778 : std_logic_vector(7 downto 0);
    signal call14_1523 : std_logic_vector(7 downto 0);
    signal call19_1535 : std_logic_vector(7 downto 0);
    signal call26_1548 : std_logic_vector(7 downto 0);
    signal call31_1560 : std_logic_vector(7 downto 0);
    signal call38_1563 : std_logic_vector(7 downto 0);
    signal call3_1498 : std_logic_vector(7 downto 0);
    signal call43_1566 : std_logic_vector(7 downto 0);
    signal call50_1580 : std_logic_vector(7 downto 0);
    signal call55_1592 : std_logic_vector(7 downto 0);
    signal call62_1605 : std_logic_vector(7 downto 0);
    signal call67_1617 : std_logic_vector(7 downto 0);
    signal call74_1620 : std_logic_vector(7 downto 0);
    signal call79_1623 : std_logic_vector(7 downto 0);
    signal call7_1510 : std_logic_vector(7 downto 0);
    signal call84_1636 : std_logic_vector(7 downto 0);
    signal call88_1648 : std_logic_vector(7 downto 0);
    signal call93_1661 : std_logic_vector(7 downto 0);
    signal call97_1673 : std_logic_vector(7 downto 0);
    signal call_1485 : std_logic_vector(7 downto 0);
    signal cmp227_1999 : std_logic_vector(0 downto 0);
    signal cmp238_2024 : std_logic_vector(0 downto 0);
    signal cmp_1969 : std_logic_vector(0 downto 0);
    signal conv102_1690 : std_logic_vector(31 downto 0);
    signal conv107_1708 : std_logic_vector(31 downto 0);
    signal conv112_1726 : std_logic_vector(31 downto 0);
    signal conv12_1514 : std_logic_vector(31 downto 0);
    signal conv131_1744 : std_logic_vector(63 downto 0);
    signal conv134_1757 : std_logic_vector(63 downto 0);
    signal conv143_1769 : std_logic_vector(63 downto 0);
    signal conv146_1782 : std_logic_vector(63 downto 0);
    signal conv15_1527 : std_logic_vector(31 downto 0);
    signal conv187_1882 : std_logic_vector(63 downto 0);
    signal conv192_1886 : std_logic_vector(63 downto 0);
    signal conv197_1890 : std_logic_vector(63 downto 0);
    signal conv211_1958 : std_logic_vector(31 downto 0);
    signal conv223_1994 : std_logic_vector(31 downto 0);
    signal conv233_2019 : std_logic_vector(31 downto 0);
    signal conv24_1539 : std_logic_vector(31 downto 0);
    signal conv27_1552 : std_logic_vector(31 downto 0);
    signal conv2_1489 : std_logic_vector(31 downto 0);
    signal conv48_1571 : std_logic_vector(15 downto 0);
    signal conv4_1502 : std_logic_vector(31 downto 0);
    signal conv51_1584 : std_logic_vector(15 downto 0);
    signal conv60_1596 : std_logic_vector(15 downto 0);
    signal conv63_1609 : std_logic_vector(15 downto 0);
    signal conv82_1627 : std_logic_vector(15 downto 0);
    signal conv85_1640 : std_logic_vector(15 downto 0);
    signal conv91_1652 : std_logic_vector(15 downto 0);
    signal conv94_1665 : std_logic_vector(15 downto 0);
    signal conv98_1677 : std_logic_vector(31 downto 0);
    signal idxprom207_1943 : std_logic_vector(63 downto 0);
    signal idxprom_1920 : std_logic_vector(63 downto 0);
    signal inc231_2003 : std_logic_vector(15 downto 0);
    signal inc231x_xinput_dim0x_x2_2008 : std_logic_vector(15 downto 0);
    signal inc_1990 : std_logic_vector(15 downto 0);
    signal indvar_1819 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2057 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2045 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1840 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2039 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1833 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2015 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2032 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1826 : std_logic_vector(15 downto 0);
    signal mul176_1873 : std_logic_vector(15 downto 0);
    signal mul198_1895 : std_logic_vector(63 downto 0);
    signal mul200_1905 : std_logic_vector(63 downto 0);
    signal mul_1863 : std_logic_vector(15 downto 0);
    signal ptr_deref_1930_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1930_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1930_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1930_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1930_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1952_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1952_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1952_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1952_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1952_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1952_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl100_1683 : std_logic_vector(31 downto 0);
    signal shl105_1701 : std_logic_vector(31 downto 0);
    signal shl110_1719 : std_logic_vector(31 downto 0);
    signal shl132_1750 : std_logic_vector(63 downto 0);
    signal shl13_1520 : std_logic_vector(31 downto 0);
    signal shl144_1775 : std_logic_vector(63 downto 0);
    signal shl25_1545 : std_logic_vector(31 downto 0);
    signal shl49_1577 : std_logic_vector(15 downto 0);
    signal shl61_1602 : std_logic_vector(15 downto 0);
    signal shl83_1633 : std_logic_vector(15 downto 0);
    signal shl92_1658 : std_logic_vector(15 downto 0);
    signal shl_1495 : std_logic_vector(31 downto 0);
    signal shr206_1937 : std_logic_vector(63 downto 0);
    signal shr237252_1816 : std_logic_vector(31 downto 0);
    signal shr_1916 : std_logic_vector(31 downto 0);
    signal sub170_1868 : std_logic_vector(15 downto 0);
    signal sub183_1810 : std_logic_vector(15 downto 0);
    signal sub184_1878 : std_logic_vector(15 downto 0);
    signal sub_1799 : std_logic_vector(15 downto 0);
    signal tmp1_1853 : std_logic_vector(31 downto 0);
    signal tmp204_1931 : std_logic_vector(63 downto 0);
    signal type_cast_1493_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1518_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1543_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1575_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1600_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1631_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1656_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1681_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1699_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1717_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1748_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1792_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1803_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1814_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1823_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1825_wire : std_logic_vector(31 downto 0);
    signal type_cast_1830_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1832_wire : std_logic_vector(15 downto 0);
    signal type_cast_1837_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1839_wire : std_logic_vector(15 downto 0);
    signal type_cast_1844_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1846_wire : std_logic_vector(15 downto 0);
    signal type_cast_1851_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1914_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1935_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1941_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1962_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1980_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1988_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2012_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2035_wire : std_logic_vector(15 downto 0);
    signal type_cast_2038_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2042_wire : std_logic_vector(15 downto 0);
    signal type_cast_2044_wire : std_logic_vector(15 downto 0);
    signal type_cast_2048_wire : std_logic_vector(15 downto 0);
    signal type_cast_2050_wire : std_logic_vector(15 downto 0);
    signal type_cast_2055_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2063_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1925_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1925_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1925_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1925_resized_base_address <= "00000000000000";
    array_obj_ref_1948_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1948_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1948_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1948_resized_base_address <= "00000000000000";
    ptr_deref_1930_word_offset_0 <= "00000000000000";
    ptr_deref_1952_word_offset_0 <= "00000000000000";
    type_cast_1493_wire_constant <= "00000000000000000000000000001000";
    type_cast_1518_wire_constant <= "00000000000000000000000000001000";
    type_cast_1543_wire_constant <= "00000000000000000000000000001000";
    type_cast_1575_wire_constant <= "0000000000001000";
    type_cast_1600_wire_constant <= "0000000000001000";
    type_cast_1631_wire_constant <= "0000000000001000";
    type_cast_1656_wire_constant <= "0000000000001000";
    type_cast_1681_wire_constant <= "00000000000000000000000000001000";
    type_cast_1699_wire_constant <= "00000000000000000000000000001000";
    type_cast_1717_wire_constant <= "00000000000000000000000000001000";
    type_cast_1748_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1792_wire_constant <= "1111111111111111";
    type_cast_1803_wire_constant <= "1111111111111111";
    type_cast_1814_wire_constant <= "00000000000000000000000000000010";
    type_cast_1823_wire_constant <= "00000000000000000000000000000000";
    type_cast_1830_wire_constant <= "0000000000000000";
    type_cast_1837_wire_constant <= "0000000000000000";
    type_cast_1844_wire_constant <= "0000000000000000";
    type_cast_1851_wire_constant <= "00000000000000000000000000000100";
    type_cast_1914_wire_constant <= "00000000000000000000000000000010";
    type_cast_1935_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1941_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1962_wire_constant <= "00000000000000000000000000000100";
    type_cast_1980_wire_constant <= "0000000000000100";
    type_cast_1988_wire_constant <= "0000000000000001";
    type_cast_2012_wire_constant <= "0000000000000000";
    type_cast_2038_wire_constant <= "0000000000000000";
    type_cast_2055_wire_constant <= "00000000000000000000000000000001";
    type_cast_2063_wire_constant <= "00000001";
    phi_stmt_1819: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1823_wire_constant & type_cast_1825_wire;
      req <= phi_stmt_1819_req_0 & phi_stmt_1819_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1819",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1819_ack_0,
          idata => idata,
          odata => indvar_1819,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1819
    phi_stmt_1826: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1830_wire_constant & type_cast_1832_wire;
      req <= phi_stmt_1826_req_0 & phi_stmt_1826_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1826",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1826_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1826,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1826
    phi_stmt_1833: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1837_wire_constant & type_cast_1839_wire;
      req <= phi_stmt_1833_req_0 & phi_stmt_1833_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1833",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1833_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1833,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1833
    phi_stmt_1840: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1844_wire_constant & type_cast_1846_wire;
      req <= phi_stmt_1840_req_0 & phi_stmt_1840_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1840",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1840_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1840,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1840
    phi_stmt_2032: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2035_wire & type_cast_2038_wire_constant;
      req <= phi_stmt_2032_req_0 & phi_stmt_2032_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2032",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2032_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2032,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2032
    phi_stmt_2039: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2042_wire & type_cast_2044_wire;
      req <= phi_stmt_2039_req_0 & phi_stmt_2039_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2039",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2039_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2039,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2039
    phi_stmt_2045: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2048_wire & type_cast_2050_wire;
      req <= phi_stmt_2045_req_0 & phi_stmt_2045_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2045",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2045_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2045,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2045
    -- flow-through select operator MUX_2014_inst
    input_dim1x_x2_2015 <= type_cast_2012_wire_constant when (cmp227_1999(0) /=  '0') else inc_1990;
    addr_of_1926_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1926_final_reg_req_0;
      addr_of_1926_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1926_final_reg_req_1;
      addr_of_1926_final_reg_ack_1<= rack(0);
      addr_of_1926_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1926_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1925_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx203_1927,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1949_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1949_final_reg_req_0;
      addr_of_1949_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1949_final_reg_req_1;
      addr_of_1949_final_reg_ack_1<= rack(0);
      addr_of_1949_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1949_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1948_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx208_1950,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1488_inst_req_0;
      type_cast_1488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1488_inst_req_1;
      type_cast_1488_inst_ack_1<= rack(0);
      type_cast_1488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_1489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1501_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1501_inst_req_0;
      type_cast_1501_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1501_inst_req_1;
      type_cast_1501_inst_ack_1<= rack(0);
      type_cast_1501_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1501_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_1502,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1513_inst_req_0;
      type_cast_1513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1513_inst_req_1;
      type_cast_1513_inst_ack_1<= rack(0);
      type_cast_1513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_1510,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1526_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1526_inst_req_0;
      type_cast_1526_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1526_inst_req_1;
      type_cast_1526_inst_ack_1<= rack(0);
      type_cast_1526_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1526_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_1523,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_1527,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1538_inst_req_0;
      type_cast_1538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1538_inst_req_1;
      type_cast_1538_inst_ack_1<= rack(0);
      type_cast_1538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_1535,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_1539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1551_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1551_inst_req_0;
      type_cast_1551_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1551_inst_req_1;
      type_cast_1551_inst_ack_1<= rack(0);
      type_cast_1551_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1551_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_1548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_1552,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1570_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1570_inst_req_0;
      type_cast_1570_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1570_inst_req_1;
      type_cast_1570_inst_ack_1<= rack(0);
      type_cast_1570_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1570_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call43_1566,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_1571,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1583_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1583_inst_req_0;
      type_cast_1583_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1583_inst_req_1;
      type_cast_1583_inst_ack_1<= rack(0);
      type_cast_1583_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1583_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_1580,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_1584,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1595_inst_req_0;
      type_cast_1595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1595_inst_req_1;
      type_cast_1595_inst_ack_1<= rack(0);
      type_cast_1595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_1592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_1596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1608_inst_req_0;
      type_cast_1608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1608_inst_req_1;
      type_cast_1608_inst_ack_1<= rack(0);
      type_cast_1608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call62_1605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_1609,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1626_inst_req_0;
      type_cast_1626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1626_inst_req_1;
      type_cast_1626_inst_ack_1<= rack(0);
      type_cast_1626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call79_1623,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_1627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1639_inst_req_0;
      type_cast_1639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1639_inst_req_1;
      type_cast_1639_inst_ack_1<= rack(0);
      type_cast_1639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call84_1636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1651_inst_req_0;
      type_cast_1651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1651_inst_req_1;
      type_cast_1651_inst_ack_1<= rack(0);
      type_cast_1651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1651_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_1648,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_1652,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1664_inst_req_0;
      type_cast_1664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1664_inst_req_1;
      type_cast_1664_inst_ack_1<= rack(0);
      type_cast_1664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_1661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1676_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1676_inst_req_0;
      type_cast_1676_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1676_inst_req_1;
      type_cast_1676_inst_ack_1<= rack(0);
      type_cast_1676_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1676_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_1673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_1677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1689_inst_req_0;
      type_cast_1689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1689_inst_req_1;
      type_cast_1689_inst_ack_1<= rack(0);
      type_cast_1689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_1686,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv102_1690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1707_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1707_inst_req_0;
      type_cast_1707_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1707_inst_req_1;
      type_cast_1707_inst_ack_1<= rack(0);
      type_cast_1707_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1707_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_1704,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1708,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1725_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1725_inst_req_0;
      type_cast_1725_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1725_inst_req_1;
      type_cast_1725_inst_ack_1<= rack(0);
      type_cast_1725_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1725_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_1722,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_1726,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1743_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1743_inst_req_0;
      type_cast_1743_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1743_inst_req_1;
      type_cast_1743_inst_ack_1<= rack(0);
      type_cast_1743_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1743_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call126_1740,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_1744,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1756_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1756_inst_req_0;
      type_cast_1756_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1756_inst_req_1;
      type_cast_1756_inst_ack_1<= rack(0);
      type_cast_1756_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1756_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_1753,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_1757,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1768_inst_req_0;
      type_cast_1768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1768_inst_req_1;
      type_cast_1768_inst_ack_1<= rack(0);
      type_cast_1768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call138_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_1769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1781_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1781_inst_req_0;
      type_cast_1781_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1781_inst_req_1;
      type_cast_1781_inst_ack_1<= rack(0);
      type_cast_1781_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1781_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_1778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv146_1782,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1825_inst_req_0;
      type_cast_1825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1825_inst_req_1;
      type_cast_1825_inst_ack_1<= rack(0);
      type_cast_1825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2057,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1825_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1832_inst_req_0;
      type_cast_1832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1832_inst_req_1;
      type_cast_1832_inst_ack_1<= rack(0);
      type_cast_1832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1832_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1839_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1839_inst_req_0;
      type_cast_1839_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1839_inst_req_1;
      type_cast_1839_inst_ack_1<= rack(0);
      type_cast_1839_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1839_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1839_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1846_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1846_inst_req_0;
      type_cast_1846_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1846_inst_req_1;
      type_cast_1846_inst_ack_1<= rack(0);
      type_cast_1846_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1846_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2045,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1846_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1881_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1881_inst_req_0;
      type_cast_1881_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1881_inst_req_1;
      type_cast_1881_inst_ack_1<= rack(0);
      type_cast_1881_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1881_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1826,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv187_1882,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1885_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1885_inst_req_0;
      type_cast_1885_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1885_inst_req_1;
      type_cast_1885_inst_ack_1<= rack(0);
      type_cast_1885_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1885_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub184_1878,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv192_1886,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1889_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1889_inst_req_0;
      type_cast_1889_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1889_inst_req_1;
      type_cast_1889_inst_ack_1<= rack(0);
      type_cast_1889_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1889_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub170_1868,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv197_1890,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1919_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1919_inst_req_0;
      type_cast_1919_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1919_inst_req_1;
      type_cast_1919_inst_ack_1<= rack(0);
      type_cast_1919_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1919_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1916,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1920,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1957_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1957_inst_req_0;
      type_cast_1957_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1957_inst_req_1;
      type_cast_1957_inst_ack_1<= rack(0);
      type_cast_1957_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1957_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1826,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_1958,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1993_inst_req_0;
      type_cast_1993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1993_inst_req_1;
      type_cast_1993_inst_ack_1<= rack(0);
      type_cast_1993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_1994,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2002_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2002_inst_req_0;
      type_cast_2002_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2002_inst_req_1;
      type_cast_2002_inst_ack_1<= rack(0);
      type_cast_2002_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2002_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp227_1999,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc231_2003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2018_inst_req_0;
      type_cast_2018_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2018_inst_req_1;
      type_cast_2018_inst_ack_1<= rack(0);
      type_cast_2018_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc231x_xinput_dim0x_x2_2008,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv233_2019,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2035_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2035_inst_req_0;
      type_cast_2035_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2035_inst_req_1;
      type_cast_2035_inst_ack_1<= rack(0);
      type_cast_2035_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2035_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add219_1982,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2035_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2042_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2042_inst_req_0;
      type_cast_2042_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2042_inst_req_1;
      type_cast_2042_inst_ack_1<= rack(0);
      type_cast_2042_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2042_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1833,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2042_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2044_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2044_inst_req_0;
      type_cast_2044_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2044_inst_req_1;
      type_cast_2044_inst_ack_1<= rack(0);
      type_cast_2044_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2044_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2015,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2044_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2048_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2048_inst_req_0;
      type_cast_2048_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2048_inst_req_1;
      type_cast_2048_inst_ack_1<= rack(0);
      type_cast_2048_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2048_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc231x_xinput_dim0x_x2_2008,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2048_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2050_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2050_inst_req_0;
      type_cast_2050_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2050_inst_req_1;
      type_cast_2050_inst_ack_1<= rack(0);
      type_cast_2050_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2050_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1840,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2050_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1925_index_1_rename
    process(R_idxprom_1924_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1924_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1924_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1925_index_1_resize
    process(idxprom_1920) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1920;
      ov := iv(13 downto 0);
      R_idxprom_1924_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1925_root_address_inst
    process(array_obj_ref_1925_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1925_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1925_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1948_index_1_rename
    process(R_idxprom207_1947_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom207_1947_resized;
      ov(13 downto 0) := iv;
      R_idxprom207_1947_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1948_index_1_resize
    process(idxprom207_1943) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom207_1943;
      ov := iv(13 downto 0);
      R_idxprom207_1947_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1948_root_address_inst
    process(array_obj_ref_1948_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1948_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1948_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1930_addr_0
    process(ptr_deref_1930_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1930_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1930_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1930_base_resize
    process(arrayidx203_1927) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx203_1927;
      ov := iv(13 downto 0);
      ptr_deref_1930_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1930_gather_scatter
    process(ptr_deref_1930_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1930_data_0;
      ov(63 downto 0) := iv;
      tmp204_1931 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1930_root_address_inst
    process(ptr_deref_1930_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1930_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1930_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1952_addr_0
    process(ptr_deref_1952_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1952_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1952_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1952_base_resize
    process(arrayidx208_1950) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx208_1950;
      ov := iv(13 downto 0);
      ptr_deref_1952_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1952_gather_scatter
    process(tmp204_1931) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp204_1931;
      ov(63 downto 0) := iv;
      ptr_deref_1952_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1952_root_address_inst
    process(ptr_deref_1952_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1952_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1952_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1970_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1969;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1970_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1970_branch_req_0,
          ack0 => if_stmt_1970_branch_ack_0,
          ack1 => if_stmt_1970_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2025_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp238_2024;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2025_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2025_branch_req_0,
          ack0 => if_stmt_2025_branch_ack_0,
          ack1 => if_stmt_2025_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1793_inst
    process(add52_1589) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add52_1589, type_cast_1792_wire_constant, tmp_var);
      add167_1794 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1804_inst
    process(add64_1614) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add64_1614, type_cast_1803_wire_constant, tmp_var);
      add180_1805 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1867_inst
    process(sub_1799, mul_1863) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1799, mul_1863, tmp_var);
      sub170_1868 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1877_inst
    process(sub183_1810, mul176_1873) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub183_1810, mul176_1873, tmp_var);
      sub184_1878 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1981_inst
    process(input_dim2x_x1_1826) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1826, type_cast_1980_wire_constant, tmp_var);
      add219_1982 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1989_inst
    process(input_dim1x_x1_1833) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1833, type_cast_1988_wire_constant, tmp_var);
      inc_1990 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2007_inst
    process(inc231_2003, input_dim0x_x2_1840) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc231_2003, input_dim0x_x2_1840, tmp_var);
      inc231x_xinput_dim0x_x2_2008 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1857_inst
    process(add113_1731, tmp1_1853) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add113_1731, tmp1_1853, tmp_var);
      add_src_0x_x0_1858 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1963_inst
    process(conv211_1958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv211_1958, type_cast_1962_wire_constant, tmp_var);
      add212_1964 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2056_inst
    process(indvar_1819) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1819, type_cast_2055_wire_constant, tmp_var);
      indvarx_xnext_2057 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1899_inst
    process(mul198_1895, conv192_1886) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul198_1895, conv192_1886, tmp_var);
      add199_1900 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1909_inst
    process(mul200_1905, conv187_1882) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul200_1905, conv187_1882, tmp_var);
      add201_1910 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1942_inst
    process(shr206_1937) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr206_1937, type_cast_1941_wire_constant, tmp_var);
      idxprom207_1943 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1998_inst
    process(conv223_1994, add16_1532) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv223_1994, add16_1532, tmp_var);
      cmp227_1999 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2023_inst
    process(conv233_2019, shr237252_1816) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv233_2019, shr237252_1816, tmp_var);
      cmp238_2024 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1815_inst
    process(add_1507) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_1507, type_cast_1814_wire_constant, tmp_var);
      shr237252_1816 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1915_inst
    process(add_src_0x_x0_1858) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1858, type_cast_1914_wire_constant, tmp_var);
      shr_1916 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1936_inst
    process(add201_1910) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add201_1910, type_cast_1935_wire_constant, tmp_var);
      shr206_1937 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1862_inst
    process(input_dim0x_x2_1840, add86_1645) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1840, add86_1645, tmp_var);
      mul_1863 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1872_inst
    process(input_dim1x_x1_1833, add86_1645) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1833, add86_1645, tmp_var);
      mul176_1873 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1852_inst
    process(indvar_1819) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1819, type_cast_1851_wire_constant, tmp_var);
      tmp1_1853 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1894_inst
    process(conv197_1890, add135_1762) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv197_1890, add135_1762, tmp_var);
      mul198_1895 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1904_inst
    process(add199_1900, add147_1787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add199_1900, add147_1787, tmp_var);
      mul200_1905 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1588_inst
    process(shl49_1577, conv51_1584) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl49_1577, conv51_1584, tmp_var);
      add52_1589 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1613_inst
    process(shl61_1602, conv63_1609) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl61_1602, conv63_1609, tmp_var);
      add64_1614 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1644_inst
    process(shl83_1633, conv85_1640) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl83_1633, conv85_1640, tmp_var);
      add86_1645 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1669_inst
    process(shl92_1658, conv94_1665) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_1658, conv94_1665, tmp_var);
      add95_1670 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1506_inst
    process(shl_1495, conv4_1502) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1495, conv4_1502, tmp_var);
      add_1507 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1531_inst
    process(shl13_1520, conv15_1527) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl13_1520, conv15_1527, tmp_var);
      add16_1532 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1556_inst
    process(shl25_1545, conv27_1552) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl25_1545, conv27_1552, tmp_var);
      add28_1557 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1694_inst
    process(shl100_1683, conv102_1690) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_1683, conv102_1690, tmp_var);
      add103_1695 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1712_inst
    process(shl105_1701, conv107_1708) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_1701, conv107_1708, tmp_var);
      add108_1713 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1730_inst
    process(shl110_1719, conv112_1726) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_1719, conv112_1726, tmp_var);
      add113_1731 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1761_inst
    process(shl132_1750, conv134_1757) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_1750, conv134_1757, tmp_var);
      add135_1762 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1786_inst
    process(shl144_1775, conv146_1782) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_1775, conv146_1782, tmp_var);
      add147_1787 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1576_inst
    process(conv48_1571) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_1571, type_cast_1575_wire_constant, tmp_var);
      shl49_1577 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1601_inst
    process(conv60_1596) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv60_1596, type_cast_1600_wire_constant, tmp_var);
      shl61_1602 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1632_inst
    process(conv82_1627) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv82_1627, type_cast_1631_wire_constant, tmp_var);
      shl83_1633 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1657_inst
    process(conv91_1652) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_1652, type_cast_1656_wire_constant, tmp_var);
      shl92_1658 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1494_inst
    process(conv2_1489) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv2_1489, type_cast_1493_wire_constant, tmp_var);
      shl_1495 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1519_inst
    process(conv12_1514) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv12_1514, type_cast_1518_wire_constant, tmp_var);
      shl13_1520 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1544_inst
    process(conv24_1539) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv24_1539, type_cast_1543_wire_constant, tmp_var);
      shl25_1545 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1682_inst
    process(conv98_1677) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv98_1677, type_cast_1681_wire_constant, tmp_var);
      shl100_1683 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1700_inst
    process(add103_1695) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add103_1695, type_cast_1699_wire_constant, tmp_var);
      shl105_1701 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1718_inst
    process(add108_1713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_1713, type_cast_1717_wire_constant, tmp_var);
      shl110_1719 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1749_inst
    process(conv131_1744) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_1744, type_cast_1748_wire_constant, tmp_var);
      shl132_1750 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1774_inst
    process(conv143_1769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv143_1769, type_cast_1773_wire_constant, tmp_var);
      shl144_1775 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1798_inst
    process(add167_1794, add95_1670) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add167_1794, add95_1670, tmp_var);
      sub_1799 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1809_inst
    process(add180_1805, add95_1670) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add180_1805, add95_1670, tmp_var);
      sub183_1810 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1968_inst
    process(add212_1964, add28_1557) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add212_1964, add28_1557, tmp_var);
      cmp_1969 <= tmp_var; --
    end process;
    -- shared split operator group (50) : array_obj_ref_1925_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1924_scaled;
      array_obj_ref_1925_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1925_index_offset_req_0;
      array_obj_ref_1925_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1925_index_offset_req_1;
      array_obj_ref_1925_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : array_obj_ref_1948_index_offset 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom207_1947_scaled;
      array_obj_ref_1948_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1948_index_offset_req_0;
      array_obj_ref_1948_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1948_index_offset_req_1;
      array_obj_ref_1948_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared load operator group (0) : ptr_deref_1930_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1930_load_0_req_0;
      ptr_deref_1930_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1930_load_0_req_1;
      ptr_deref_1930_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1930_word_address_0;
      ptr_deref_1930_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1952_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1952_store_0_req_0;
      ptr_deref_1952_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1952_store_0_req_1;
      ptr_deref_1952_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1952_word_address_0;
      data_in <= ptr_deref_1952_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1562_inst RPIPE_Block0_start_1522_inst RPIPE_Block0_start_1604_inst RPIPE_Block0_start_1685_inst RPIPE_Block0_start_1559_inst RPIPE_Block0_start_1509_inst RPIPE_Block0_start_1591_inst RPIPE_Block0_start_1660_inst RPIPE_Block0_start_1622_inst RPIPE_Block0_start_1497_inst RPIPE_Block0_start_1484_inst RPIPE_Block0_start_1619_inst RPIPE_Block0_start_1547_inst RPIPE_Block0_start_1635_inst RPIPE_Block0_start_1647_inst RPIPE_Block0_start_1616_inst RPIPE_Block0_start_1534_inst RPIPE_Block0_start_1672_inst RPIPE_Block0_start_1565_inst RPIPE_Block0_start_1579_inst RPIPE_Block0_start_1703_inst RPIPE_Block0_start_1721_inst RPIPE_Block0_start_1733_inst RPIPE_Block0_start_1736_inst RPIPE_Block0_start_1739_inst RPIPE_Block0_start_1752_inst RPIPE_Block0_start_1764_inst RPIPE_Block0_start_1777_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 27 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 27 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant outBUFs : IntegerArray(27 downto 0) := (27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      reqL_unguarded(27) <= RPIPE_Block0_start_1562_inst_req_0;
      reqL_unguarded(26) <= RPIPE_Block0_start_1522_inst_req_0;
      reqL_unguarded(25) <= RPIPE_Block0_start_1604_inst_req_0;
      reqL_unguarded(24) <= RPIPE_Block0_start_1685_inst_req_0;
      reqL_unguarded(23) <= RPIPE_Block0_start_1559_inst_req_0;
      reqL_unguarded(22) <= RPIPE_Block0_start_1509_inst_req_0;
      reqL_unguarded(21) <= RPIPE_Block0_start_1591_inst_req_0;
      reqL_unguarded(20) <= RPIPE_Block0_start_1660_inst_req_0;
      reqL_unguarded(19) <= RPIPE_Block0_start_1622_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Block0_start_1497_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Block0_start_1484_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Block0_start_1619_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Block0_start_1547_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Block0_start_1635_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Block0_start_1647_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1616_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1534_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1672_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1565_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1579_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1703_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1721_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1733_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1736_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1739_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1752_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1764_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1777_inst_req_0;
      RPIPE_Block0_start_1562_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_Block0_start_1522_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_Block0_start_1604_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_Block0_start_1685_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_Block0_start_1559_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_Block0_start_1509_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_Block0_start_1591_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_Block0_start_1660_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_Block0_start_1622_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Block0_start_1497_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Block0_start_1484_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Block0_start_1619_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Block0_start_1547_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Block0_start_1635_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Block0_start_1647_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1616_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1534_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1672_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1565_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1579_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1703_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1721_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1733_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1736_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1739_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1752_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1764_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1777_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(27) <= RPIPE_Block0_start_1562_inst_req_1;
      reqR_unguarded(26) <= RPIPE_Block0_start_1522_inst_req_1;
      reqR_unguarded(25) <= RPIPE_Block0_start_1604_inst_req_1;
      reqR_unguarded(24) <= RPIPE_Block0_start_1685_inst_req_1;
      reqR_unguarded(23) <= RPIPE_Block0_start_1559_inst_req_1;
      reqR_unguarded(22) <= RPIPE_Block0_start_1509_inst_req_1;
      reqR_unguarded(21) <= RPIPE_Block0_start_1591_inst_req_1;
      reqR_unguarded(20) <= RPIPE_Block0_start_1660_inst_req_1;
      reqR_unguarded(19) <= RPIPE_Block0_start_1622_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Block0_start_1497_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Block0_start_1484_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Block0_start_1619_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Block0_start_1547_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Block0_start_1635_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Block0_start_1647_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1616_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1534_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1672_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1565_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1579_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1703_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1721_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1733_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1736_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1739_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1752_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1764_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1777_inst_req_1;
      RPIPE_Block0_start_1562_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_Block0_start_1522_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_Block0_start_1604_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_Block0_start_1685_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_Block0_start_1559_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_Block0_start_1509_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_Block0_start_1591_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_Block0_start_1660_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_Block0_start_1622_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Block0_start_1497_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Block0_start_1484_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Block0_start_1619_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Block0_start_1547_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Block0_start_1635_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Block0_start_1647_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1616_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1534_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1672_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1565_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1579_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1703_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1721_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1733_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1736_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1739_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1752_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1764_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1777_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      call38_1563 <= data_out(223 downto 216);
      call14_1523 <= data_out(215 downto 208);
      call62_1605 <= data_out(207 downto 200);
      call101_1686 <= data_out(199 downto 192);
      call31_1560 <= data_out(191 downto 184);
      call7_1510 <= data_out(183 downto 176);
      call55_1592 <= data_out(175 downto 168);
      call93_1661 <= data_out(167 downto 160);
      call79_1623 <= data_out(159 downto 152);
      call3_1498 <= data_out(151 downto 144);
      call_1485 <= data_out(143 downto 136);
      call74_1620 <= data_out(135 downto 128);
      call26_1548 <= data_out(127 downto 120);
      call84_1636 <= data_out(119 downto 112);
      call88_1648 <= data_out(111 downto 104);
      call67_1617 <= data_out(103 downto 96);
      call19_1535 <= data_out(95 downto 88);
      call97_1673 <= data_out(87 downto 80);
      call43_1566 <= data_out(79 downto 72);
      call50_1580 <= data_out(71 downto 64);
      call106_1704 <= data_out(63 downto 56);
      call111_1722 <= data_out(55 downto 48);
      call114_1734 <= data_out(47 downto 40);
      call121_1737 <= data_out(39 downto 32);
      call126_1740 <= data_out(31 downto 24);
      call133_1753 <= data_out(23 downto 16);
      call138_1765 <= data_out(15 downto 8);
      call145_1778 <= data_out(7 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 8,  num_reqs => 28,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_2061_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_2061_inst_req_0;
      WPIPE_Block0_done_2061_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_2061_inst_req_1;
      WPIPE_Block0_done_2061_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2063_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_5537_start: Boolean;
  signal convTransposeB_CP_5537_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_2272_inst_req_0 : boolean;
  signal type_cast_2276_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2290_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2272_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2320_inst_ack_1 : boolean;
  signal type_cast_2276_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2326_inst_ack_0 : boolean;
  signal type_cast_2330_inst_ack_0 : boolean;
  signal type_cast_2263_inst_ack_1 : boolean;
  signal type_cast_2343_inst_req_0 : boolean;
  signal type_cast_2263_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2320_inst_req_1 : boolean;
  signal type_cast_2330_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2364_inst_ack_0 : boolean;
  signal type_cast_2294_inst_req_0 : boolean;
  signal type_cast_2294_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2326_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2290_inst_ack_1 : boolean;
  signal type_cast_2312_inst_req_0 : boolean;
  signal type_cast_2312_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2320_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2351_inst_req_1 : boolean;
  signal type_cast_2312_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2320_inst_req_0 : boolean;
  signal type_cast_2312_inst_req_1 : boolean;
  signal type_cast_2481_inst_ack_1 : boolean;
  signal type_cast_2477_inst_req_0 : boolean;
  signal type_cast_2477_inst_ack_0 : boolean;
  signal type_cast_2294_inst_req_1 : boolean;
  signal type_cast_2485_inst_req_1 : boolean;
  signal type_cast_2485_inst_ack_1 : boolean;
  signal type_cast_2276_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2326_inst_req_1 : boolean;
  signal type_cast_2276_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2351_inst_req_0 : boolean;
  signal type_cast_2368_inst_ack_0 : boolean;
  signal type_cast_2294_inst_ack_1 : boolean;
  signal type_cast_2406_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2339_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2290_inst_ack_0 : boolean;
  signal type_cast_2355_inst_req_1 : boolean;
  signal type_cast_2355_inst_ack_1 : boolean;
  signal type_cast_2368_inst_req_1 : boolean;
  signal type_cast_2406_inst_req_0 : boolean;
  signal type_cast_2481_inst_req_0 : boolean;
  signal type_cast_2481_inst_ack_0 : boolean;
  signal type_cast_2406_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2272_inst_ack_1 : boolean;
  signal type_cast_2481_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2339_inst_ack_0 : boolean;
  signal type_cast_2343_inst_ack_0 : boolean;
  signal type_cast_2368_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2272_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2351_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2308_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2308_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2326_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2351_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2323_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2364_inst_req_1 : boolean;
  signal type_cast_2485_inst_req_0 : boolean;
  signal type_cast_2485_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2364_inst_ack_1 : boolean;
  signal type_cast_2368_inst_req_0 : boolean;
  signal type_cast_2330_inst_req_1 : boolean;
  signal type_cast_2355_inst_req_0 : boolean;
  signal type_cast_2355_inst_ack_0 : boolean;
  signal type_cast_2330_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2364_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2290_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2308_inst_req_1 : boolean;
  signal type_cast_2477_inst_req_1 : boolean;
  signal type_cast_2477_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2308_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2323_inst_req_0 : boolean;
  signal type_cast_2406_inst_ack_0 : boolean;
  signal type_cast_2343_inst_req_1 : boolean;
  signal type_cast_2343_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2323_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2339_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2339_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2323_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2072_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2072_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2072_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2072_inst_ack_1 : boolean;
  signal type_cast_2076_inst_req_0 : boolean;
  signal type_cast_2076_inst_ack_0 : boolean;
  signal type_cast_2076_inst_req_1 : boolean;
  signal type_cast_2076_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2085_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2085_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2085_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2085_inst_ack_1 : boolean;
  signal type_cast_2089_inst_req_0 : boolean;
  signal type_cast_2089_inst_ack_0 : boolean;
  signal type_cast_2089_inst_req_1 : boolean;
  signal type_cast_2089_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2097_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2097_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2097_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2097_inst_ack_1 : boolean;
  signal type_cast_2101_inst_req_0 : boolean;
  signal type_cast_2101_inst_ack_0 : boolean;
  signal type_cast_2101_inst_req_1 : boolean;
  signal type_cast_2101_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2110_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2110_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2110_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2110_inst_ack_1 : boolean;
  signal type_cast_2114_inst_req_0 : boolean;
  signal type_cast_2114_inst_ack_0 : boolean;
  signal type_cast_2114_inst_req_1 : boolean;
  signal type_cast_2114_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2122_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2122_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2122_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2122_inst_ack_1 : boolean;
  signal type_cast_2126_inst_req_0 : boolean;
  signal type_cast_2126_inst_ack_0 : boolean;
  signal type_cast_2126_inst_req_1 : boolean;
  signal type_cast_2126_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2135_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2135_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2135_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2135_inst_ack_1 : boolean;
  signal type_cast_2139_inst_req_0 : boolean;
  signal type_cast_2139_inst_ack_0 : boolean;
  signal type_cast_2139_inst_req_1 : boolean;
  signal type_cast_2139_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2147_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2147_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2147_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2147_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2150_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2150_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2150_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2150_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2153_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2153_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2153_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2153_inst_ack_1 : boolean;
  signal type_cast_2157_inst_req_0 : boolean;
  signal type_cast_2157_inst_ack_0 : boolean;
  signal type_cast_2157_inst_req_1 : boolean;
  signal type_cast_2157_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2166_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2166_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2166_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2166_inst_ack_1 : boolean;
  signal type_cast_2170_inst_req_0 : boolean;
  signal type_cast_2170_inst_ack_0 : boolean;
  signal type_cast_2170_inst_req_1 : boolean;
  signal type_cast_2170_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2178_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2178_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2178_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2178_inst_ack_1 : boolean;
  signal type_cast_2182_inst_req_0 : boolean;
  signal type_cast_2182_inst_ack_0 : boolean;
  signal type_cast_2182_inst_req_1 : boolean;
  signal type_cast_2182_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2191_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2191_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2191_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2191_inst_ack_1 : boolean;
  signal type_cast_2195_inst_req_0 : boolean;
  signal type_cast_2195_inst_ack_0 : boolean;
  signal type_cast_2195_inst_req_1 : boolean;
  signal type_cast_2195_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2203_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2203_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2203_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2203_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2206_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2206_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2206_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2206_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2209_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2209_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2209_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2209_inst_ack_1 : boolean;
  signal type_cast_2213_inst_req_0 : boolean;
  signal type_cast_2213_inst_ack_0 : boolean;
  signal type_cast_2213_inst_req_1 : boolean;
  signal type_cast_2213_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2222_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2222_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2222_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2222_inst_ack_1 : boolean;
  signal type_cast_2226_inst_req_0 : boolean;
  signal type_cast_2226_inst_ack_0 : boolean;
  signal type_cast_2226_inst_req_1 : boolean;
  signal type_cast_2226_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2234_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2234_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2234_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2234_inst_ack_1 : boolean;
  signal type_cast_2238_inst_req_0 : boolean;
  signal type_cast_2238_inst_ack_0 : boolean;
  signal type_cast_2238_inst_req_1 : boolean;
  signal type_cast_2238_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2247_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2247_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2247_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2247_inst_ack_1 : boolean;
  signal type_cast_2251_inst_req_0 : boolean;
  signal type_cast_2251_inst_ack_0 : boolean;
  signal type_cast_2251_inst_req_1 : boolean;
  signal type_cast_2251_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_2259_inst_req_0 : boolean;
  signal RPIPE_Block1_start_2259_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_2259_inst_req_1 : boolean;
  signal RPIPE_Block1_start_2259_inst_ack_1 : boolean;
  signal type_cast_2263_inst_req_0 : boolean;
  signal type_cast_2263_inst_ack_0 : boolean;
  signal type_cast_2515_inst_req_0 : boolean;
  signal type_cast_2515_inst_ack_0 : boolean;
  signal type_cast_2515_inst_req_1 : boolean;
  signal type_cast_2515_inst_ack_1 : boolean;
  signal array_obj_ref_2521_index_offset_req_0 : boolean;
  signal array_obj_ref_2521_index_offset_ack_0 : boolean;
  signal array_obj_ref_2521_index_offset_req_1 : boolean;
  signal array_obj_ref_2521_index_offset_ack_1 : boolean;
  signal addr_of_2522_final_reg_req_0 : boolean;
  signal addr_of_2522_final_reg_ack_0 : boolean;
  signal addr_of_2522_final_reg_req_1 : boolean;
  signal addr_of_2522_final_reg_ack_1 : boolean;
  signal ptr_deref_2526_load_0_req_0 : boolean;
  signal ptr_deref_2526_load_0_ack_0 : boolean;
  signal ptr_deref_2526_load_0_req_1 : boolean;
  signal ptr_deref_2526_load_0_ack_1 : boolean;
  signal array_obj_ref_2544_index_offset_req_0 : boolean;
  signal array_obj_ref_2544_index_offset_ack_0 : boolean;
  signal array_obj_ref_2544_index_offset_req_1 : boolean;
  signal array_obj_ref_2544_index_offset_ack_1 : boolean;
  signal addr_of_2545_final_reg_req_0 : boolean;
  signal addr_of_2545_final_reg_ack_0 : boolean;
  signal addr_of_2545_final_reg_req_1 : boolean;
  signal addr_of_2545_final_reg_ack_1 : boolean;
  signal ptr_deref_2548_store_0_req_0 : boolean;
  signal ptr_deref_2548_store_0_ack_0 : boolean;
  signal ptr_deref_2548_store_0_req_1 : boolean;
  signal ptr_deref_2548_store_0_ack_1 : boolean;
  signal type_cast_2553_inst_req_0 : boolean;
  signal type_cast_2553_inst_ack_0 : boolean;
  signal type_cast_2553_inst_req_1 : boolean;
  signal type_cast_2553_inst_ack_1 : boolean;
  signal if_stmt_2566_branch_req_0 : boolean;
  signal if_stmt_2566_branch_ack_1 : boolean;
  signal if_stmt_2566_branch_ack_0 : boolean;
  signal type_cast_2589_inst_req_0 : boolean;
  signal type_cast_2589_inst_ack_0 : boolean;
  signal type_cast_2589_inst_req_1 : boolean;
  signal type_cast_2589_inst_ack_1 : boolean;
  signal type_cast_2598_inst_req_0 : boolean;
  signal type_cast_2598_inst_ack_0 : boolean;
  signal type_cast_2598_inst_req_1 : boolean;
  signal type_cast_2598_inst_ack_1 : boolean;
  signal type_cast_2614_inst_req_0 : boolean;
  signal type_cast_2614_inst_ack_0 : boolean;
  signal type_cast_2614_inst_req_1 : boolean;
  signal type_cast_2614_inst_ack_1 : boolean;
  signal if_stmt_2621_branch_req_0 : boolean;
  signal if_stmt_2621_branch_ack_1 : boolean;
  signal if_stmt_2621_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2657_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2657_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2657_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2657_inst_ack_1 : boolean;
  signal phi_stmt_2416_req_0 : boolean;
  signal phi_stmt_2423_req_1 : boolean;
  signal phi_stmt_2430_req_1 : boolean;
  signal type_cast_2442_inst_req_0 : boolean;
  signal type_cast_2442_inst_ack_0 : boolean;
  signal type_cast_2442_inst_req_1 : boolean;
  signal type_cast_2442_inst_ack_1 : boolean;
  signal phi_stmt_2437_req_1 : boolean;
  signal type_cast_2422_inst_req_0 : boolean;
  signal type_cast_2422_inst_ack_0 : boolean;
  signal type_cast_2422_inst_req_1 : boolean;
  signal type_cast_2422_inst_ack_1 : boolean;
  signal phi_stmt_2416_req_1 : boolean;
  signal type_cast_2426_inst_req_0 : boolean;
  signal type_cast_2426_inst_ack_0 : boolean;
  signal type_cast_2426_inst_req_1 : boolean;
  signal type_cast_2426_inst_ack_1 : boolean;
  signal phi_stmt_2423_req_0 : boolean;
  signal type_cast_2433_inst_req_0 : boolean;
  signal type_cast_2433_inst_ack_0 : boolean;
  signal type_cast_2433_inst_req_1 : boolean;
  signal type_cast_2433_inst_ack_1 : boolean;
  signal phi_stmt_2430_req_0 : boolean;
  signal type_cast_2440_inst_req_0 : boolean;
  signal type_cast_2440_inst_ack_0 : boolean;
  signal type_cast_2440_inst_req_1 : boolean;
  signal type_cast_2440_inst_ack_1 : boolean;
  signal phi_stmt_2437_req_0 : boolean;
  signal phi_stmt_2416_ack_0 : boolean;
  signal phi_stmt_2423_ack_0 : boolean;
  signal phi_stmt_2430_ack_0 : boolean;
  signal phi_stmt_2437_ack_0 : boolean;
  signal phi_stmt_2628_req_0 : boolean;
  signal type_cast_2638_inst_req_0 : boolean;
  signal type_cast_2638_inst_ack_0 : boolean;
  signal type_cast_2638_inst_req_1 : boolean;
  signal type_cast_2638_inst_ack_1 : boolean;
  signal phi_stmt_2635_req_0 : boolean;
  signal type_cast_2644_inst_req_0 : boolean;
  signal type_cast_2644_inst_ack_0 : boolean;
  signal type_cast_2644_inst_req_1 : boolean;
  signal type_cast_2644_inst_ack_1 : boolean;
  signal phi_stmt_2641_req_0 : boolean;
  signal type_cast_2634_inst_req_0 : boolean;
  signal type_cast_2634_inst_ack_0 : boolean;
  signal type_cast_2634_inst_req_1 : boolean;
  signal type_cast_2634_inst_ack_1 : boolean;
  signal phi_stmt_2628_req_1 : boolean;
  signal type_cast_2640_inst_req_0 : boolean;
  signal type_cast_2640_inst_ack_0 : boolean;
  signal type_cast_2640_inst_req_1 : boolean;
  signal type_cast_2640_inst_ack_1 : boolean;
  signal phi_stmt_2635_req_1 : boolean;
  signal type_cast_2646_inst_req_0 : boolean;
  signal type_cast_2646_inst_ack_0 : boolean;
  signal type_cast_2646_inst_req_1 : boolean;
  signal type_cast_2646_inst_ack_1 : boolean;
  signal phi_stmt_2641_req_1 : boolean;
  signal phi_stmt_2628_ack_0 : boolean;
  signal phi_stmt_2635_ack_0 : boolean;
  signal phi_stmt_2641_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_5537_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5537_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_5537_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5537_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_5537: Block -- control-path 
    signal convTransposeB_CP_5537_elements: BooleanArray(190 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_5537_elements(0) <= convTransposeB_CP_5537_start;
    convTransposeB_CP_5537_symbol <= convTransposeB_CP_5537_elements(141);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0:  members (74) 
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2070/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/branch_block_stmt_2070__entry__
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_update_start_
      -- 
    cr_6052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2263_inst_req_1); -- 
    cr_6136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2312_inst_req_1); -- 
    cr_6108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2294_inst_req_1); -- 
    cr_6080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2276_inst_req_1); -- 
    cr_6248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2355_inst_req_1); -- 
    cr_6276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2368_inst_req_1); -- 
    cr_6192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2330_inst_req_1); -- 
    cr_6220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2343_inst_req_1); -- 
    rr_5585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => RPIPE_Block1_start_2072_inst_req_0); -- 
    cr_5604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2076_inst_req_1); -- 
    cr_5632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2089_inst_req_1); -- 
    cr_5660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2101_inst_req_1); -- 
    cr_5688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2114_inst_req_1); -- 
    cr_5716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2126_inst_req_1); -- 
    cr_5744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2139_inst_req_1); -- 
    cr_5800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2157_inst_req_1); -- 
    cr_5828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2170_inst_req_1); -- 
    cr_5856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2182_inst_req_1); -- 
    cr_5884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2195_inst_req_1); -- 
    cr_5940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2213_inst_req_1); -- 
    cr_5968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2226_inst_req_1); -- 
    cr_5996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2238_inst_req_1); -- 
    cr_6024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(0), ack => type_cast_2251_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	190 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	155 
    -- CP-element group 1: 	149 
    -- CP-element group 1: 	150 
    -- CP-element group 1: 	159 
    -- CP-element group 1: 	156 
    -- CP-element group 1: 	153 
    -- CP-element group 1: 	158 
    -- CP-element group 1: 	152 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2070/merge_stmt_2627__exit__
      -- CP-element group 1: 	 branch_block_stmt_2070/assign_stmt_2653__entry__
      -- CP-element group 1: 	 branch_block_stmt_2070/assign_stmt_2653__exit__
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2070/assign_stmt_2653/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/assign_stmt_2653/$exit
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/Update/cr
      -- 
    rr_6734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(1), ack => type_cast_2422_inst_req_0); -- 
    cr_6739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(1), ack => type_cast_2422_inst_req_1); -- 
    rr_6757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(1), ack => type_cast_2426_inst_req_0); -- 
    cr_6762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(1), ack => type_cast_2426_inst_req_1); -- 
    rr_6780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(1), ack => type_cast_2433_inst_req_0); -- 
    cr_6785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(1), ack => type_cast_2433_inst_req_1); -- 
    rr_6803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(1), ack => type_cast_2440_inst_req_0); -- 
    cr_6808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(1), ack => type_cast_2440_inst_req_1); -- 
    convTransposeB_CP_5537_elements(1) <= convTransposeB_CP_5537_elements(190);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_Update/cr
      -- 
    ra_5586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2072_inst_ack_0, ack => convTransposeB_CP_5537_elements(2)); -- 
    cr_5590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(2), ack => RPIPE_Block1_start_2072_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2072_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_Sample/rr
      -- 
    ca_5591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2072_inst_ack_1, ack => convTransposeB_CP_5537_elements(3)); -- 
    rr_5599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(3), ack => type_cast_2076_inst_req_0); -- 
    rr_5613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(3), ack => RPIPE_Block1_start_2085_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_Sample/ra
      -- 
    ra_5600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2076_inst_ack_0, ack => convTransposeB_CP_5537_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	102 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2076_Update/ca
      -- 
    ca_5605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2076_inst_ack_1, ack => convTransposeB_CP_5537_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_Update/cr
      -- 
    ra_5614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2085_inst_ack_0, ack => convTransposeB_CP_5537_elements(6)); -- 
    cr_5618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(6), ack => RPIPE_Block1_start_2085_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2085_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_Sample/rr
      -- 
    ca_5619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2085_inst_ack_1, ack => convTransposeB_CP_5537_elements(7)); -- 
    rr_5627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(7), ack => type_cast_2089_inst_req_0); -- 
    rr_5641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(7), ack => RPIPE_Block1_start_2097_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_Sample/ra
      -- 
    ra_5628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2089_inst_ack_0, ack => convTransposeB_CP_5537_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	102 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2089_Update/ca
      -- 
    ca_5633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2089_inst_ack_1, ack => convTransposeB_CP_5537_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_Update/cr
      -- 
    ra_5642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2097_inst_ack_0, ack => convTransposeB_CP_5537_elements(10)); -- 
    cr_5646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(10), ack => RPIPE_Block1_start_2097_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2097_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_Sample/rr
      -- 
    ca_5647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2097_inst_ack_1, ack => convTransposeB_CP_5537_elements(11)); -- 
    rr_5655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(11), ack => type_cast_2101_inst_req_0); -- 
    rr_5669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(11), ack => RPIPE_Block1_start_2110_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_Sample/ra
      -- 
    ra_5656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2101_inst_ack_0, ack => convTransposeB_CP_5537_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	102 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2101_Update/ca
      -- 
    ca_5661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2101_inst_ack_1, ack => convTransposeB_CP_5537_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_Update/cr
      -- 
    ra_5670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2110_inst_ack_0, ack => convTransposeB_CP_5537_elements(14)); -- 
    cr_5674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(14), ack => RPIPE_Block1_start_2110_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2110_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_Sample/rr
      -- 
    ca_5675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2110_inst_ack_1, ack => convTransposeB_CP_5537_elements(15)); -- 
    rr_5683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(15), ack => type_cast_2114_inst_req_0); -- 
    rr_5697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(15), ack => RPIPE_Block1_start_2122_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_Sample/ra
      -- 
    ra_5684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2114_inst_ack_0, ack => convTransposeB_CP_5537_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	102 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2114_Update/ca
      -- 
    ca_5689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2114_inst_ack_1, ack => convTransposeB_CP_5537_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_Update/cr
      -- 
    ra_5698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2122_inst_ack_0, ack => convTransposeB_CP_5537_elements(18)); -- 
    cr_5702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(18), ack => RPIPE_Block1_start_2122_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2122_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_Sample/rr
      -- 
    ca_5703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2122_inst_ack_1, ack => convTransposeB_CP_5537_elements(19)); -- 
    rr_5711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(19), ack => type_cast_2126_inst_req_0); -- 
    rr_5725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(19), ack => RPIPE_Block1_start_2135_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_Sample/ra
      -- 
    ra_5712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2126_inst_ack_0, ack => convTransposeB_CP_5537_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	102 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2126_Update/ca
      -- 
    ca_5717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2126_inst_ack_1, ack => convTransposeB_CP_5537_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_update_start_
      -- CP-element group 22: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_Update/cr
      -- 
    ra_5726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2135_inst_ack_0, ack => convTransposeB_CP_5537_elements(22)); -- 
    cr_5730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(22), ack => RPIPE_Block1_start_2135_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2135_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_Sample/rr
      -- 
    ca_5731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2135_inst_ack_1, ack => convTransposeB_CP_5537_elements(23)); -- 
    rr_5739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(23), ack => type_cast_2139_inst_req_0); -- 
    rr_5753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(23), ack => RPIPE_Block1_start_2147_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_Sample/ra
      -- 
    ra_5740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2139_inst_ack_0, ack => convTransposeB_CP_5537_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	102 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2139_Update/ca
      -- 
    ca_5745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2139_inst_ack_1, ack => convTransposeB_CP_5537_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_update_start_
      -- CP-element group 26: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_Update/cr
      -- 
    ra_5754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2147_inst_ack_0, ack => convTransposeB_CP_5537_elements(26)); -- 
    cr_5758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(26), ack => RPIPE_Block1_start_2147_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2147_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_Sample/rr
      -- 
    ca_5759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2147_inst_ack_1, ack => convTransposeB_CP_5537_elements(27)); -- 
    rr_5767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(27), ack => RPIPE_Block1_start_2150_inst_req_0); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_Update/cr
      -- 
    ra_5768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2150_inst_ack_0, ack => convTransposeB_CP_5537_elements(28)); -- 
    cr_5772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(28), ack => RPIPE_Block1_start_2150_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2150_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_Sample/rr
      -- 
    ca_5773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2150_inst_ack_1, ack => convTransposeB_CP_5537_elements(29)); -- 
    rr_5781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(29), ack => RPIPE_Block1_start_2153_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_Update/cr
      -- 
    ra_5782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2153_inst_ack_0, ack => convTransposeB_CP_5537_elements(30)); -- 
    cr_5786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(30), ack => RPIPE_Block1_start_2153_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2153_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_Sample/rr
      -- 
    ca_5787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2153_inst_ack_1, ack => convTransposeB_CP_5537_elements(31)); -- 
    rr_5809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(31), ack => RPIPE_Block1_start_2166_inst_req_0); -- 
    rr_5795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(31), ack => type_cast_2157_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_Sample/ra
      -- 
    ra_5796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2157_inst_ack_0, ack => convTransposeB_CP_5537_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	102 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2157_Update/ca
      -- 
    ca_5801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2157_inst_ack_1, ack => convTransposeB_CP_5537_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_Update/cr
      -- 
    ra_5810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2166_inst_ack_0, ack => convTransposeB_CP_5537_elements(34)); -- 
    cr_5814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(34), ack => RPIPE_Block1_start_2166_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2166_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_Sample/rr
      -- 
    ca_5815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2166_inst_ack_1, ack => convTransposeB_CP_5537_elements(35)); -- 
    rr_5823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(35), ack => type_cast_2170_inst_req_0); -- 
    rr_5837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(35), ack => RPIPE_Block1_start_2178_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_Sample/ra
      -- 
    ra_5824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2170_inst_ack_0, ack => convTransposeB_CP_5537_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	102 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2170_Update/ca
      -- 
    ca_5829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2170_inst_ack_1, ack => convTransposeB_CP_5537_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_update_start_
      -- CP-element group 38: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_Update/cr
      -- 
    ra_5838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2178_inst_ack_0, ack => convTransposeB_CP_5537_elements(38)); -- 
    cr_5842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(38), ack => RPIPE_Block1_start_2178_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	42 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2178_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_Sample/rr
      -- 
    ca_5843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2178_inst_ack_1, ack => convTransposeB_CP_5537_elements(39)); -- 
    rr_5865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(39), ack => RPIPE_Block1_start_2191_inst_req_0); -- 
    rr_5851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(39), ack => type_cast_2182_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_Sample/ra
      -- 
    ra_5852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2182_inst_ack_0, ack => convTransposeB_CP_5537_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	102 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2182_Update/ca
      -- 
    ca_5857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2182_inst_ack_1, ack => convTransposeB_CP_5537_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_update_start_
      -- CP-element group 42: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_Update/cr
      -- 
    ra_5866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2191_inst_ack_0, ack => convTransposeB_CP_5537_elements(42)); -- 
    cr_5870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(42), ack => RPIPE_Block1_start_2191_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	46 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2191_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_Sample/rr
      -- 
    ca_5871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2191_inst_ack_1, ack => convTransposeB_CP_5537_elements(43)); -- 
    rr_5893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(43), ack => RPIPE_Block1_start_2203_inst_req_0); -- 
    rr_5879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(43), ack => type_cast_2195_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_Sample/ra
      -- 
    ra_5880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2195_inst_ack_0, ack => convTransposeB_CP_5537_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	102 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2195_Update/ca
      -- 
    ca_5885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2195_inst_ack_1, ack => convTransposeB_CP_5537_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_update_start_
      -- CP-element group 46: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_Update/cr
      -- 
    ra_5894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2203_inst_ack_0, ack => convTransposeB_CP_5537_elements(46)); -- 
    cr_5898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(46), ack => RPIPE_Block1_start_2203_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2203_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_Sample/rr
      -- 
    ca_5899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2203_inst_ack_1, ack => convTransposeB_CP_5537_elements(47)); -- 
    rr_5907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(47), ack => RPIPE_Block1_start_2206_inst_req_0); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_update_start_
      -- CP-element group 48: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_Update/cr
      -- 
    ra_5908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2206_inst_ack_0, ack => convTransposeB_CP_5537_elements(48)); -- 
    cr_5912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(48), ack => RPIPE_Block1_start_2206_inst_req_1); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2206_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_Sample/rr
      -- 
    ca_5913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2206_inst_ack_1, ack => convTransposeB_CP_5537_elements(49)); -- 
    rr_5921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(49), ack => RPIPE_Block1_start_2209_inst_req_0); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_update_start_
      -- CP-element group 50: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_Update/cr
      -- 
    ra_5922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2209_inst_ack_0, ack => convTransposeB_CP_5537_elements(50)); -- 
    cr_5926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(50), ack => RPIPE_Block1_start_2209_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2209_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_Sample/rr
      -- 
    ca_5927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2209_inst_ack_1, ack => convTransposeB_CP_5537_elements(51)); -- 
    rr_5949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(51), ack => RPIPE_Block1_start_2222_inst_req_0); -- 
    rr_5935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(51), ack => type_cast_2213_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_Sample/ra
      -- 
    ra_5936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2213_inst_ack_0, ack => convTransposeB_CP_5537_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	102 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2213_Update/ca
      -- 
    ca_5941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2213_inst_ack_1, ack => convTransposeB_CP_5537_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_update_start_
      -- CP-element group 54: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_Update/cr
      -- 
    ra_5950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2222_inst_ack_0, ack => convTransposeB_CP_5537_elements(54)); -- 
    cr_5954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(54), ack => RPIPE_Block1_start_2222_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2222_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_Sample/rr
      -- 
    ca_5955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2222_inst_ack_1, ack => convTransposeB_CP_5537_elements(55)); -- 
    rr_5977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(55), ack => RPIPE_Block1_start_2234_inst_req_0); -- 
    rr_5963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(55), ack => type_cast_2226_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_Sample/ra
      -- 
    ra_5964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2226_inst_ack_0, ack => convTransposeB_CP_5537_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	102 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2226_Update/ca
      -- 
    ca_5969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2226_inst_ack_1, ack => convTransposeB_CP_5537_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_update_start_
      -- CP-element group 58: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_Update/cr
      -- 
    ra_5978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2234_inst_ack_0, ack => convTransposeB_CP_5537_elements(58)); -- 
    cr_5982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(58), ack => RPIPE_Block1_start_2234_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2234_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_Sample/rr
      -- 
    ca_5983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2234_inst_ack_1, ack => convTransposeB_CP_5537_elements(59)); -- 
    rr_6005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(59), ack => RPIPE_Block1_start_2247_inst_req_0); -- 
    rr_5991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(59), ack => type_cast_2238_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_Sample/ra
      -- 
    ra_5992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2238_inst_ack_0, ack => convTransposeB_CP_5537_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	102 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2238_Update/ca
      -- 
    ca_5997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2238_inst_ack_1, ack => convTransposeB_CP_5537_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_Update/cr
      -- 
    ra_6006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2247_inst_ack_0, ack => convTransposeB_CP_5537_elements(62)); -- 
    cr_6010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(62), ack => RPIPE_Block1_start_2247_inst_req_1); -- 
    -- CP-element group 63:  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2247_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_Sample/rr
      -- 
    ca_6011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2247_inst_ack_1, ack => convTransposeB_CP_5537_elements(63)); -- 
    rr_6019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(63), ack => type_cast_2251_inst_req_0); -- 
    rr_6033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(63), ack => RPIPE_Block1_start_2259_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_Sample/ra
      -- 
    ra_6020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2251_inst_ack_0, ack => convTransposeB_CP_5537_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	102 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2251_Update/ca
      -- 
    ca_6025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2251_inst_ack_1, ack => convTransposeB_CP_5537_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_update_start_
      -- CP-element group 66: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_Update/cr
      -- 
    ra_6034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2259_inst_ack_0, ack => convTransposeB_CP_5537_elements(66)); -- 
    cr_6038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(66), ack => RPIPE_Block1_start_2259_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2259_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_Sample/rr
      -- 
    ca_6039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2259_inst_ack_1, ack => convTransposeB_CP_5537_elements(67)); -- 
    rr_6047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(67), ack => type_cast_2263_inst_req_0); -- 
    rr_6061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(67), ack => RPIPE_Block1_start_2272_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_Sample/ra
      -- 
    ra_6048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2263_inst_ack_0, ack => convTransposeB_CP_5537_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	102 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_Update/ca
      -- CP-element group 69: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2263_update_completed_
      -- 
    ca_6053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2263_inst_ack_1, ack => convTransposeB_CP_5537_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_Update/$entry
      -- 
    ra_6062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2272_inst_ack_0, ack => convTransposeB_CP_5537_elements(70)); -- 
    cr_6066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(70), ack => RPIPE_Block1_start_2272_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	74 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2272_Update/$exit
      -- 
    ca_6067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2272_inst_ack_1, ack => convTransposeB_CP_5537_elements(71)); -- 
    rr_6075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(71), ack => type_cast_2276_inst_req_0); -- 
    rr_6089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(71), ack => RPIPE_Block1_start_2290_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_sample_completed_
      -- 
    ra_6076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2276_inst_ack_0, ack => convTransposeB_CP_5537_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	102 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2276_update_completed_
      -- 
    ca_6081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2276_inst_ack_1, ack => convTransposeB_CP_5537_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	71 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_Update/cr
      -- CP-element group 74: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_update_start_
      -- 
    ra_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2290_inst_ack_0, ack => convTransposeB_CP_5537_elements(74)); -- 
    cr_6094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(74), ack => RPIPE_Block1_start_2290_inst_req_1); -- 
    -- CP-element group 75:  fork  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (9) 
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2290_Update/$exit
      -- 
    ca_6095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2290_inst_ack_1, ack => convTransposeB_CP_5537_elements(75)); -- 
    rr_6117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(75), ack => RPIPE_Block1_start_2308_inst_req_0); -- 
    rr_6103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(75), ack => type_cast_2294_inst_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_Sample/ra
      -- 
    ra_6104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2294_inst_ack_0, ack => convTransposeB_CP_5537_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	102 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2294_Update/ca
      -- 
    ca_6109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2294_inst_ack_1, ack => convTransposeB_CP_5537_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_Update/cr
      -- 
    ra_6118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2308_inst_ack_0, ack => convTransposeB_CP_5537_elements(78)); -- 
    cr_6122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(78), ack => RPIPE_Block1_start_2308_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2308_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_Sample/$entry
      -- 
    ca_6123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2308_inst_ack_1, ack => convTransposeB_CP_5537_elements(79)); -- 
    rr_6145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(79), ack => RPIPE_Block1_start_2320_inst_req_0); -- 
    rr_6131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(79), ack => type_cast_2312_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_Sample/$exit
      -- 
    ra_6132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_0, ack => convTransposeB_CP_5537_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	102 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2312_Update/$exit
      -- 
    ca_6137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_1, ack => convTransposeB_CP_5537_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_update_start_
      -- CP-element group 82: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_Sample/ra
      -- 
    ra_6146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2320_inst_ack_0, ack => convTransposeB_CP_5537_elements(82)); -- 
    cr_6150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(82), ack => RPIPE_Block1_start_2320_inst_req_1); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2320_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_Sample/rr
      -- 
    ca_6151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2320_inst_ack_1, ack => convTransposeB_CP_5537_elements(83)); -- 
    rr_6159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(83), ack => RPIPE_Block1_start_2323_inst_req_0); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_update_start_
      -- CP-element group 84: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_Update/cr
      -- 
    ra_6160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2323_inst_ack_0, ack => convTransposeB_CP_5537_elements(84)); -- 
    cr_6164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(84), ack => RPIPE_Block1_start_2323_inst_req_1); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2323_Update/ca
      -- 
    ca_6165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2323_inst_ack_1, ack => convTransposeB_CP_5537_elements(85)); -- 
    rr_6173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(85), ack => RPIPE_Block1_start_2326_inst_req_0); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_sample_completed_
      -- 
    ra_6174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2326_inst_ack_0, ack => convTransposeB_CP_5537_elements(86)); -- 
    cr_6178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(86), ack => RPIPE_Block1_start_2326_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	90 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2326_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_sample_start_
      -- 
    ca_6179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2326_inst_ack_1, ack => convTransposeB_CP_5537_elements(87)); -- 
    rr_6201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(87), ack => RPIPE_Block1_start_2339_inst_req_0); -- 
    rr_6187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(87), ack => type_cast_2330_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_sample_completed_
      -- 
    ra_6188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2330_inst_ack_0, ack => convTransposeB_CP_5537_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	102 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2330_Update/ca
      -- 
    ca_6193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2330_inst_ack_1, ack => convTransposeB_CP_5537_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_update_start_
      -- CP-element group 90: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_Update/cr
      -- 
    ra_6202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2339_inst_ack_0, ack => convTransposeB_CP_5537_elements(90)); -- 
    cr_6206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(90), ack => RPIPE_Block1_start_2339_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	94 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2339_Update/ca
      -- 
    ca_6207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2339_inst_ack_1, ack => convTransposeB_CP_5537_elements(91)); -- 
    rr_6229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(91), ack => RPIPE_Block1_start_2351_inst_req_0); -- 
    rr_6215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(91), ack => type_cast_2343_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_Sample/ra
      -- 
    ra_6216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2343_inst_ack_0, ack => convTransposeB_CP_5537_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	102 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2343_Update/ca
      -- 
    ca_6221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2343_inst_ack_1, ack => convTransposeB_CP_5537_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_update_start_
      -- CP-element group 94: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_Update/$entry
      -- 
    ra_6230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2351_inst_ack_0, ack => convTransposeB_CP_5537_elements(94)); -- 
    cr_6234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(94), ack => RPIPE_Block1_start_2351_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2351_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_Sample/rr
      -- 
    ca_6235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2351_inst_ack_1, ack => convTransposeB_CP_5537_elements(95)); -- 
    rr_6257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(95), ack => RPIPE_Block1_start_2364_inst_req_0); -- 
    rr_6243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(95), ack => type_cast_2355_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_Sample/ra
      -- 
    ra_6244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2355_inst_ack_0, ack => convTransposeB_CP_5537_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	102 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2355_update_completed_
      -- 
    ca_6249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2355_inst_ack_1, ack => convTransposeB_CP_5537_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_Update/$entry
      -- 
    ra_6258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2364_inst_ack_0, ack => convTransposeB_CP_5537_elements(98)); -- 
    cr_6262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(98), ack => RPIPE_Block1_start_2364_inst_req_1); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/RPIPE_Block1_start_2364_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_sample_start_
      -- 
    ca_6263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_2364_inst_ack_1, ack => convTransposeB_CP_5537_elements(99)); -- 
    rr_6271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(99), ack => type_cast_2368_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_Sample/$exit
      -- 
    ra_6272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2368_inst_ack_0, ack => convTransposeB_CP_5537_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/type_cast_2368_update_completed_
      -- 
    ca_6277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2368_inst_ack_1, ack => convTransposeB_CP_5537_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	101 
    -- CP-element group 102: 	77 
    -- CP-element group 102: 	33 
    -- CP-element group 102: 	89 
    -- CP-element group 102: 	97 
    -- CP-element group 102: 	93 
    -- CP-element group 102: 	81 
    -- CP-element group 102: 	73 
    -- CP-element group 102: 	69 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	61 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	41 
    -- CP-element group 102: 	37 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	5 
    -- CP-element group 102: 	9 
    -- CP-element group 102: 	13 
    -- CP-element group 102: 	17 
    -- CP-element group 102: 	21 
    -- CP-element group 102: 	25 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (10) 
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413__entry__
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374__exit__
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/$entry
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_update_start_
      -- CP-element group 102: 	 branch_block_stmt_2070/assign_stmt_2073_to_assign_stmt_2374/$exit
      -- 
    rr_6288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(102), ack => type_cast_2406_inst_req_0); -- 
    cr_6293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(102), ack => type_cast_2406_inst_req_1); -- 
    convTransposeB_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(65) & convTransposeB_CP_5537_elements(101) & convTransposeB_CP_5537_elements(77) & convTransposeB_CP_5537_elements(33) & convTransposeB_CP_5537_elements(89) & convTransposeB_CP_5537_elements(97) & convTransposeB_CP_5537_elements(93) & convTransposeB_CP_5537_elements(81) & convTransposeB_CP_5537_elements(73) & convTransposeB_CP_5537_elements(69) & convTransposeB_CP_5537_elements(53) & convTransposeB_CP_5537_elements(61) & convTransposeB_CP_5537_elements(45) & convTransposeB_CP_5537_elements(41) & convTransposeB_CP_5537_elements(37) & convTransposeB_CP_5537_elements(57) & convTransposeB_CP_5537_elements(5) & convTransposeB_CP_5537_elements(9) & convTransposeB_CP_5537_elements(13) & convTransposeB_CP_5537_elements(17) & convTransposeB_CP_5537_elements(21) & convTransposeB_CP_5537_elements(25);
      gj_convTransposeB_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_Sample/ra
      -- 
    ra_6289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2406_inst_ack_0, ack => convTransposeB_CP_5537_elements(103)); -- 
    -- CP-element group 104:  fork  transition  place  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	146 
    -- CP-element group 104: 	145 
    -- CP-element group 104: 	142 
    -- CP-element group 104: 	143 
    -- CP-element group 104: 	144 
    -- CP-element group 104:  members (21) 
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody
      -- CP-element group 104: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413__exit__
      -- CP-element group 104: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/$exit
      -- CP-element group 104: 	 branch_block_stmt_2070/assign_stmt_2381_to_assign_stmt_2413/type_cast_2406_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2416/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2423/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2430/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/Update/cr
      -- 
    ca_6294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2406_inst_ack_1, ack => convTransposeB_CP_5537_elements(104)); -- 
    rr_6708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(104), ack => type_cast_2442_inst_req_0); -- 
    cr_6713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(104), ack => type_cast_2442_inst_req_1); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	167 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_sample_completed_
      -- 
    ra_6306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2477_inst_ack_0, ack => convTransposeB_CP_5537_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	167 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	119 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_Update/ca
      -- 
    ca_6311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2477_inst_ack_1, ack => convTransposeB_CP_5537_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	167 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_Sample/$exit
      -- 
    ra_6320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2481_inst_ack_0, ack => convTransposeB_CP_5537_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	167 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_update_completed_
      -- 
    ca_6325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2481_inst_ack_1, ack => convTransposeB_CP_5537_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	167 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_Sample/$exit
      -- 
    ra_6334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2485_inst_ack_0, ack => convTransposeB_CP_5537_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	167 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	119 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_update_completed_
      -- 
    ca_6339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2485_inst_ack_1, ack => convTransposeB_CP_5537_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	167 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_Sample/ra
      -- 
    ra_6348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2515_inst_ack_0, ack => convTransposeB_CP_5537_elements(111)); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	167 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (16) 
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_resized_1
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_scaled_1
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_computed_1
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_resize_1/$entry
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_resize_1/$exit
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_resize_1/index_resize_req
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_resize_1/index_resize_ack
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_scale_1/$entry
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_scale_1/$exit
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_scale_1/scale_rename_req
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_index_scale_1/scale_rename_ack
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_Sample/req
      -- 
    ca_6353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2515_inst_ack_1, ack => convTransposeB_CP_5537_elements(112)); -- 
    req_6378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(112), ack => array_obj_ref_2521_index_offset_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	129 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_sample_complete
      -- CP-element group 113: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_Sample/ack
      -- 
    ack_6379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2521_index_offset_ack_0, ack => convTransposeB_CP_5537_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	167 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (11) 
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_root_address_calculated
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_offset_calculated
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_Update/ack
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_base_plus_offset/$entry
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_base_plus_offset/$exit
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_base_plus_offset/sum_rename_req
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_base_plus_offset/sum_rename_ack
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_request/$entry
      -- CP-element group 114: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_request/req
      -- 
    ack_6384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2521_index_offset_ack_1, ack => convTransposeB_CP_5537_elements(114)); -- 
    req_6393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(114), ack => addr_of_2522_final_reg_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_request/$exit
      -- CP-element group 115: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_request/ack
      -- 
    ack_6394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2522_final_reg_ack_0, ack => convTransposeB_CP_5537_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	167 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (24) 
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_complete/$exit
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_complete/ack
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_word_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_root_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_address_resized
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_addr_resize/$entry
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_addr_resize/$exit
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_addr_resize/base_resize_req
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_addr_resize/base_resize_ack
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_plus_offset/$entry
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_plus_offset/$exit
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_plus_offset/sum_rename_req
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_base_plus_offset/sum_rename_ack
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_word_addrgen/$entry
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_word_addrgen/$exit
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_word_addrgen/root_register_req
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_word_addrgen/root_register_ack
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Sample/word_access_start/$entry
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Sample/word_access_start/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Sample/word_access_start/word_0/rr
      -- 
    ack_6399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2522_final_reg_ack_1, ack => convTransposeB_CP_5537_elements(116)); -- 
    rr_6432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(116), ack => ptr_deref_2526_load_0_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Sample/word_access_start/word_0/ra
      -- 
    ra_6433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2526_load_0_ack_0, ack => convTransposeB_CP_5537_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	167 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	124 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/ptr_deref_2526_Merge/$entry
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/ptr_deref_2526_Merge/$exit
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/ptr_deref_2526_Merge/merge_req
      -- CP-element group 118: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/ptr_deref_2526_Merge/merge_ack
      -- 
    ca_6444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2526_load_0_ack_1, ack => convTransposeB_CP_5537_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	110 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	106 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (13) 
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_scale_1/$entry
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_resized_1
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_scaled_1
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_computed_1
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_resize_1/$entry
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_resize_1/$exit
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_resize_1/index_resize_req
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_resize_1/index_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_scale_1/$exit
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_scale_1/scale_rename_req
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_index_scale_1/scale_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_Sample/req
      -- 
    req_6474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(119), ack => array_obj_ref_2544_index_offset_req_0); -- 
    convTransposeB_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(110) & convTransposeB_CP_5537_elements(108) & convTransposeB_CP_5537_elements(106);
      gj_convTransposeB_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	129 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_sample_complete
      -- CP-element group 120: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_Sample/ack
      -- 
    ack_6475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2544_index_offset_ack_0, ack => convTransposeB_CP_5537_elements(120)); -- 
    -- CP-element group 121:  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (11) 
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_root_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_offset_calculated
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_Update/ack
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_base_plus_offset/$entry
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_base_plus_offset/$exit
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_base_plus_offset/sum_rename_req
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_base_plus_offset/sum_rename_ack
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_request/$entry
      -- CP-element group 121: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_request/req
      -- 
    ack_6480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2544_index_offset_ack_1, ack => convTransposeB_CP_5537_elements(121)); -- 
    req_6489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(121), ack => addr_of_2545_final_reg_req_0); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_request/$exit
      -- CP-element group 122: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_request/ack
      -- 
    ack_6490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2545_final_reg_ack_0, ack => convTransposeB_CP_5537_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	167 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (19) 
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_complete/$exit
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_complete/ack
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_word_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_root_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_address_resized
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_addr_resize/$entry
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_addr_resize/$exit
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_addr_resize/base_resize_req
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_addr_resize/base_resize_ack
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_plus_offset/$entry
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_plus_offset/$exit
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_plus_offset/sum_rename_req
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_base_plus_offset/sum_rename_ack
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_word_addrgen/$entry
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_word_addrgen/$exit
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_word_addrgen/root_register_req
      -- CP-element group 123: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_word_addrgen/root_register_ack
      -- 
    ack_6495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2545_final_reg_ack_1, ack => convTransposeB_CP_5537_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: 	118 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/ptr_deref_2548_Split/$entry
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/ptr_deref_2548_Split/$exit
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/ptr_deref_2548_Split/split_req
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/ptr_deref_2548_Split/split_ack
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/word_access_start/$entry
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/word_access_start/word_0/$entry
      -- CP-element group 124: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/word_access_start/word_0/rr
      -- 
    rr_6533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(124), ack => ptr_deref_2548_store_0_req_0); -- 
    convTransposeB_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(123) & convTransposeB_CP_5537_elements(118);
      gj_convTransposeB_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/word_access_start/$exit
      -- CP-element group 125: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/word_access_start/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Sample/word_access_start/word_0/ra
      -- 
    ra_6534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2548_store_0_ack_0, ack => convTransposeB_CP_5537_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	167 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	129 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Update/word_access_complete/$exit
      -- CP-element group 126: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Update/word_access_complete/word_0/$exit
      -- CP-element group 126: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Update/word_access_complete/word_0/ca
      -- 
    ca_6545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2548_store_0_ack_1, ack => convTransposeB_CP_5537_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	167 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_Sample/ra
      -- 
    ra_6554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2553_inst_ack_0, ack => convTransposeB_CP_5537_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	167 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_Update/ca
      -- 
    ca_6559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2553_inst_ack_1, ack => convTransposeB_CP_5537_elements(128)); -- 
    -- CP-element group 129:  branch  join  transition  place  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	126 
    -- CP-element group 129: 	120 
    -- CP-element group 129: 	113 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (10) 
      -- CP-element group 129: 	 branch_block_stmt_2070/if_stmt_2566__entry__
      -- CP-element group 129: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565__exit__
      -- CP-element group 129: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/$exit
      -- CP-element group 129: 	 branch_block_stmt_2070/if_stmt_2566_dead_link/$entry
      -- CP-element group 129: 	 branch_block_stmt_2070/if_stmt_2566_eval_test/$entry
      -- CP-element group 129: 	 branch_block_stmt_2070/if_stmt_2566_eval_test/$exit
      -- CP-element group 129: 	 branch_block_stmt_2070/if_stmt_2566_eval_test/branch_req
      -- CP-element group 129: 	 branch_block_stmt_2070/R_cmp_2567_place
      -- CP-element group 129: 	 branch_block_stmt_2070/if_stmt_2566_if_link/$entry
      -- CP-element group 129: 	 branch_block_stmt_2070/if_stmt_2566_else_link/$entry
      -- 
    branch_req_6567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(129), ack => if_stmt_2566_branch_req_0); -- 
    convTransposeB_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(126) & convTransposeB_CP_5537_elements(120) & convTransposeB_CP_5537_elements(113) & convTransposeB_CP_5537_elements(128);
      gj_convTransposeB_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	179 
    -- CP-element group 130: 	180 
    -- CP-element group 130: 	182 
    -- CP-element group 130: 	176 
    -- CP-element group 130: 	177 
    -- CP-element group 130: 	183 
    -- CP-element group 130:  members (40) 
      -- CP-element group 130: 	 branch_block_stmt_2070/merge_stmt_2572__exit__
      -- CP-element group 130: 	 branch_block_stmt_2070/assign_stmt_2578__entry__
      -- CP-element group 130: 	 branch_block_stmt_2070/assign_stmt_2578__exit__
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254
      -- CP-element group 130: 	 branch_block_stmt_2070/if_stmt_2566_if_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_2070/if_stmt_2566_if_link/if_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_2070/whilex_xbody_ifx_xthen
      -- CP-element group 130: 	 branch_block_stmt_2070/assign_stmt_2578/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/assign_stmt_2578/$exit
      -- CP-element group 130: 	 branch_block_stmt_2070/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_2070/merge_stmt_2572_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_2070/merge_stmt_2572_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/merge_stmt_2572_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_2070/merge_stmt_2572_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/Update/cr
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/Update/cr
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2566_branch_ack_1, ack => convTransposeB_CP_5537_elements(130)); -- 
    rr_6918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(130), ack => type_cast_2634_inst_req_0); -- 
    cr_6923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(130), ack => type_cast_2634_inst_req_1); -- 
    rr_6941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(130), ack => type_cast_2640_inst_req_0); -- 
    cr_6946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(130), ack => type_cast_2640_inst_req_1); -- 
    rr_6964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(130), ack => type_cast_2646_inst_req_0); -- 
    cr_6969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(130), ack => type_cast_2646_inst_req_1); -- 
    -- CP-element group 131:  fork  transition  place  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	137 
    -- CP-element group 131: 	135 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (24) 
      -- CP-element group 131: 	 branch_block_stmt_2070/merge_stmt_2580__exit__
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620__entry__
      -- CP-element group 131: 	 branch_block_stmt_2070/if_stmt_2566_else_link/$exit
      -- CP-element group 131: 	 branch_block_stmt_2070/if_stmt_2566_else_link/else_choice_transition
      -- CP-element group 131: 	 branch_block_stmt_2070/whilex_xbody_ifx_xelse
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/$entry
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_update_start_
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_update_start_
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_update_start_
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_2070/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 131: 	 branch_block_stmt_2070/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 131: 	 branch_block_stmt_2070/merge_stmt_2580_PhiReqMerge
      -- CP-element group 131: 	 branch_block_stmt_2070/merge_stmt_2580_PhiAck/$entry
      -- CP-element group 131: 	 branch_block_stmt_2070/merge_stmt_2580_PhiAck/$exit
      -- CP-element group 131: 	 branch_block_stmt_2070/merge_stmt_2580_PhiAck/dummy
      -- 
    else_choice_transition_6576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2566_branch_ack_0, ack => convTransposeB_CP_5537_elements(131)); -- 
    rr_6592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(131), ack => type_cast_2589_inst_req_0); -- 
    cr_6597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(131), ack => type_cast_2589_inst_req_1); -- 
    cr_6611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(131), ack => type_cast_2598_inst_req_1); -- 
    cr_6625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(131), ack => type_cast_2614_inst_req_1); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_Sample/ra
      -- 
    ra_6593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_0, ack => convTransposeB_CP_5537_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2589_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_Sample/rr
      -- 
    ca_6598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_1, ack => convTransposeB_CP_5537_elements(133)); -- 
    rr_6606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(133), ack => type_cast_2598_inst_req_0); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_Sample/ra
      -- 
    ra_6607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2598_inst_ack_0, ack => convTransposeB_CP_5537_elements(134)); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	131 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (6) 
      -- CP-element group 135: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2598_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_Sample/rr
      -- 
    ca_6612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2598_inst_ack_1, ack => convTransposeB_CP_5537_elements(135)); -- 
    rr_6620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(135), ack => type_cast_2614_inst_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_Sample/ra
      -- 
    ra_6621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_0, ack => convTransposeB_CP_5537_elements(136)); -- 
    -- CP-element group 137:  branch  transition  place  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	131 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (13) 
      -- CP-element group 137: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620__exit__
      -- CP-element group 137: 	 branch_block_stmt_2070/if_stmt_2621__entry__
      -- CP-element group 137: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/$exit
      -- CP-element group 137: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_2070/assign_stmt_2586_to_assign_stmt_2620/type_cast_2614_Update/ca
      -- CP-element group 137: 	 branch_block_stmt_2070/if_stmt_2621_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_2070/if_stmt_2621_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_2070/if_stmt_2621_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_2070/if_stmt_2621_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_2070/R_cmp243_2622_place
      -- CP-element group 137: 	 branch_block_stmt_2070/if_stmt_2621_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_2070/if_stmt_2621_else_link/$entry
      -- 
    ca_6626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2614_inst_ack_1, ack => convTransposeB_CP_5537_elements(137)); -- 
    branch_req_6634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(137), ack => if_stmt_2621_branch_req_0); -- 
    -- CP-element group 138:  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (15) 
      -- CP-element group 138: 	 branch_block_stmt_2070/merge_stmt_2655__exit__
      -- CP-element group 138: 	 branch_block_stmt_2070/assign_stmt_2660__entry__
      -- CP-element group 138: 	 branch_block_stmt_2070/if_stmt_2621_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_2070/if_stmt_2621_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_2070/ifx_xelse_whilex_xend
      -- CP-element group 138: 	 branch_block_stmt_2070/assign_stmt_2660/$entry
      -- CP-element group 138: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_Sample/req
      -- CP-element group 138: 	 branch_block_stmt_2070/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_2070/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 138: 	 branch_block_stmt_2070/merge_stmt_2655_PhiReqMerge
      -- CP-element group 138: 	 branch_block_stmt_2070/merge_stmt_2655_PhiAck/$entry
      -- CP-element group 138: 	 branch_block_stmt_2070/merge_stmt_2655_PhiAck/$exit
      -- CP-element group 138: 	 branch_block_stmt_2070/merge_stmt_2655_PhiAck/dummy
      -- 
    if_choice_transition_6639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2621_branch_ack_1, ack => convTransposeB_CP_5537_elements(138)); -- 
    req_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(138), ack => WPIPE_Block1_done_2657_inst_req_0); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	172 
    -- CP-element group 139: 	173 
    -- CP-element group 139: 	169 
    -- CP-element group 139: 	168 
    -- CP-element group 139: 	170 
    -- CP-element group 139:  members (22) 
      -- CP-element group 139: 	 branch_block_stmt_2070/if_stmt_2621_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_2070/if_stmt_2621_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2628/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/Update/cr
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2621_branch_ack_0, ack => convTransposeB_CP_5537_elements(139)); -- 
    rr_6869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(139), ack => type_cast_2638_inst_req_0); -- 
    cr_6874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(139), ack => type_cast_2638_inst_req_1); -- 
    rr_6892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(139), ack => type_cast_2644_inst_req_0); -- 
    cr_6897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(139), ack => type_cast_2644_inst_req_1); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (6) 
      -- CP-element group 140: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_update_start_
      -- CP-element group 140: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_Sample/ack
      -- CP-element group 140: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_Update/req
      -- 
    ack_6660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2657_inst_ack_0, ack => convTransposeB_CP_5537_elements(140)); -- 
    req_6664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(140), ack => WPIPE_Block1_done_2657_inst_req_1); -- 
    -- CP-element group 141:  transition  place  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (16) 
      -- CP-element group 141: 	 branch_block_stmt_2070/branch_block_stmt_2070__exit__
      -- CP-element group 141: 	 branch_block_stmt_2070/$exit
      -- CP-element group 141: 	 $exit
      -- CP-element group 141: 	 branch_block_stmt_2070/assign_stmt_2660__exit__
      -- CP-element group 141: 	 branch_block_stmt_2070/return__
      -- CP-element group 141: 	 branch_block_stmt_2070/merge_stmt_2662__exit__
      -- CP-element group 141: 	 branch_block_stmt_2070/assign_stmt_2660/$exit
      -- CP-element group 141: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_2070/assign_stmt_2660/WPIPE_Block1_done_2657_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_2070/return___PhiReq/$entry
      -- CP-element group 141: 	 branch_block_stmt_2070/return___PhiReq/$exit
      -- CP-element group 141: 	 branch_block_stmt_2070/merge_stmt_2662_PhiReqMerge
      -- CP-element group 141: 	 branch_block_stmt_2070/merge_stmt_2662_PhiAck/$entry
      -- CP-element group 141: 	 branch_block_stmt_2070/merge_stmt_2662_PhiAck/$exit
      -- CP-element group 141: 	 branch_block_stmt_2070/merge_stmt_2662_PhiAck/dummy
      -- 
    ack_6665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2657_inst_ack_1, ack => convTransposeB_CP_5537_elements(141)); -- 
    -- CP-element group 142:  transition  output  delay-element  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	104 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	148 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2416/$exit
      -- CP-element group 142: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/$exit
      -- CP-element group 142: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2420_konst_delay_trans
      -- CP-element group 142: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_req
      -- 
    phi_stmt_2416_req_6676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2416_req_6676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(142), ack => phi_stmt_2416_req_0); -- 
    -- Element group convTransposeB_CP_5537_elements(142) is a control-delay.
    cp_element_142_delay: control_delay_element  generic map(name => " 142_delay", delay_value => 1)  port map(req => convTransposeB_CP_5537_elements(104), ack => convTransposeB_CP_5537_elements(142), clk => clk, reset =>reset);
    -- CP-element group 143:  transition  output  delay-element  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	104 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	148 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2423/$exit
      -- CP-element group 143: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/$exit
      -- CP-element group 143: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2429_konst_delay_trans
      -- CP-element group 143: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_req
      -- 
    phi_stmt_2423_req_6684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2423_req_6684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(143), ack => phi_stmt_2423_req_1); -- 
    -- Element group convTransposeB_CP_5537_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => convTransposeB_CP_5537_elements(104), ack => convTransposeB_CP_5537_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  transition  output  delay-element  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	104 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	148 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2430/$exit
      -- CP-element group 144: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/$exit
      -- CP-element group 144: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2436_konst_delay_trans
      -- CP-element group 144: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_req
      -- 
    phi_stmt_2430_req_6692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2430_req_6692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(144), ack => phi_stmt_2430_req_1); -- 
    -- Element group convTransposeB_CP_5537_elements(144) is a control-delay.
    cp_element_144_delay: control_delay_element  generic map(name => " 144_delay", delay_value => 1)  port map(req => convTransposeB_CP_5537_elements(104), ack => convTransposeB_CP_5537_elements(144), clk => clk, reset =>reset);
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	104 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/Sample/ra
      -- 
    ra_6709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2442_inst_ack_0, ack => convTransposeB_CP_5537_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	104 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/Update/ca
      -- 
    ca_6714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2442_inst_ack_1, ack => convTransposeB_CP_5537_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/$exit
      -- CP-element group 147: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/$exit
      -- CP-element group 147: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/$exit
      -- CP-element group 147: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2442/SplitProtocol/$exit
      -- CP-element group 147: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_req
      -- 
    phi_stmt_2437_req_6715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2437_req_6715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(147), ack => phi_stmt_2437_req_1); -- 
    convTransposeB_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(146) & convTransposeB_CP_5537_elements(145);
      gj_convTransposeB_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: 	142 
    -- CP-element group 148: 	143 
    -- CP-element group 148: 	144 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	162 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_2070/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(147) & convTransposeB_CP_5537_elements(142) & convTransposeB_CP_5537_elements(143) & convTransposeB_CP_5537_elements(144);
      gj_convTransposeB_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	1 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/Sample/ra
      -- 
    ra_6735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2422_inst_ack_0, ack => convTransposeB_CP_5537_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	1 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (2) 
      -- CP-element group 150: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/Update/ca
      -- 
    ca_6740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2422_inst_ack_1, ack => convTransposeB_CP_5537_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	161 
    -- CP-element group 151:  members (5) 
      -- CP-element group 151: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/$exit
      -- CP-element group 151: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/$exit
      -- CP-element group 151: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/$exit
      -- CP-element group 151: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_sources/type_cast_2422/SplitProtocol/$exit
      -- CP-element group 151: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2416/phi_stmt_2416_req
      -- 
    phi_stmt_2416_req_6741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2416_req_6741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(151), ack => phi_stmt_2416_req_1); -- 
    convTransposeB_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(149) & convTransposeB_CP_5537_elements(150);
      gj_convTransposeB_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	1 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/Sample/ra
      -- 
    ra_6758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2426_inst_ack_0, ack => convTransposeB_CP_5537_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	1 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/Update/ca
      -- 
    ca_6763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2426_inst_ack_1, ack => convTransposeB_CP_5537_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	161 
    -- CP-element group 154:  members (5) 
      -- CP-element group 154: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/$exit
      -- CP-element group 154: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/$exit
      -- CP-element group 154: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/$exit
      -- CP-element group 154: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_sources/type_cast_2426/SplitProtocol/$exit
      -- CP-element group 154: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2423/phi_stmt_2423_req
      -- 
    phi_stmt_2423_req_6764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2423_req_6764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(154), ack => phi_stmt_2423_req_0); -- 
    convTransposeB_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(153) & convTransposeB_CP_5537_elements(152);
      gj_convTransposeB_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	1 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (2) 
      -- CP-element group 155: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/Sample/ra
      -- 
    ra_6781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2433_inst_ack_0, ack => convTransposeB_CP_5537_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	1 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/Update/ca
      -- 
    ca_6786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2433_inst_ack_1, ack => convTransposeB_CP_5537_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	161 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/$exit
      -- CP-element group 157: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/$exit
      -- CP-element group 157: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/$exit
      -- CP-element group 157: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_sources/type_cast_2433/SplitProtocol/$exit
      -- CP-element group 157: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2430/phi_stmt_2430_req
      -- 
    phi_stmt_2430_req_6787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2430_req_6787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(157), ack => phi_stmt_2430_req_0); -- 
    convTransposeB_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(155) & convTransposeB_CP_5537_elements(156);
      gj_convTransposeB_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	1 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (2) 
      -- CP-element group 158: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/Sample/ra
      -- 
    ra_6804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2440_inst_ack_0, ack => convTransposeB_CP_5537_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	1 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/Update/ca
      -- 
    ca_6809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2440_inst_ack_1, ack => convTransposeB_CP_5537_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (5) 
      -- CP-element group 160: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/$exit
      -- CP-element group 160: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/$exit
      -- CP-element group 160: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/$exit
      -- CP-element group 160: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_sources/type_cast_2440/SplitProtocol/$exit
      -- CP-element group 160: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/phi_stmt_2437/phi_stmt_2437_req
      -- 
    phi_stmt_2437_req_6810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2437_req_6810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(160), ack => phi_stmt_2437_req_0); -- 
    convTransposeB_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(159) & convTransposeB_CP_5537_elements(158);
      gj_convTransposeB_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	151 
    -- CP-element group 161: 	160 
    -- CP-element group 161: 	157 
    -- CP-element group 161: 	154 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_2070/ifx_xend254_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(151) & convTransposeB_CP_5537_elements(160) & convTransposeB_CP_5537_elements(157) & convTransposeB_CP_5537_elements(154);
      gj_convTransposeB_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  merge  fork  transition  place  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	148 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	164 
    -- CP-element group 162: 	165 
    -- CP-element group 162: 	166 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_2070/merge_stmt_2415_PhiReqMerge
      -- CP-element group 162: 	 branch_block_stmt_2070/merge_stmt_2415_PhiAck/$entry
      -- 
    convTransposeB_CP_5537_elements(162) <= OrReduce(convTransposeB_CP_5537_elements(148) & convTransposeB_CP_5537_elements(161));
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	167 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_2070/merge_stmt_2415_PhiAck/phi_stmt_2416_ack
      -- 
    phi_stmt_2416_ack_6815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2416_ack_0, ack => convTransposeB_CP_5537_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	167 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_2070/merge_stmt_2415_PhiAck/phi_stmt_2423_ack
      -- 
    phi_stmt_2423_ack_6816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2423_ack_0, ack => convTransposeB_CP_5537_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	162 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (1) 
      -- CP-element group 165: 	 branch_block_stmt_2070/merge_stmt_2415_PhiAck/phi_stmt_2430_ack
      -- 
    phi_stmt_2430_ack_6817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2430_ack_0, ack => convTransposeB_CP_5537_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	162 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_2070/merge_stmt_2415_PhiAck/phi_stmt_2437_ack
      -- 
    phi_stmt_2437_ack_6818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2437_ack_0, ack => convTransposeB_CP_5537_elements(166)); -- 
    -- CP-element group 167:  join  fork  transition  place  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	163 
    -- CP-element group 167: 	164 
    -- CP-element group 167: 	165 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	123 
    -- CP-element group 167: 	116 
    -- CP-element group 167: 	112 
    -- CP-element group 167: 	110 
    -- CP-element group 167: 	107 
    -- CP-element group 167: 	108 
    -- CP-element group 167: 	126 
    -- CP-element group 167: 	111 
    -- CP-element group 167: 	118 
    -- CP-element group 167: 	127 
    -- CP-element group 167: 	121 
    -- CP-element group 167: 	128 
    -- CP-element group 167: 	114 
    -- CP-element group 167: 	105 
    -- CP-element group 167: 	106 
    -- CP-element group 167: 	109 
    -- CP-element group 167:  members (56) 
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565__entry__
      -- CP-element group 167: 	 branch_block_stmt_2070/merge_stmt_2415__exit__
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2485_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2477_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2481_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2515_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_update_start
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2521_final_index_sum_regn_Update/req
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2522_complete/req
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/word_access_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/word_access_complete/word_0/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2526_Update/word_access_complete/word_0/cr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_update_start
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/array_obj_ref_2544_final_index_sum_regn_Update/req
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/addr_of_2545_complete/req
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Update/word_access_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Update/word_access_complete/word_0/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/ptr_deref_2548_Update/word_access_complete/word_0/cr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2070/assign_stmt_2449_to_assign_stmt_2565/type_cast_2553_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2070/merge_stmt_2415_PhiAck/$exit
      -- 
    rr_6305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2477_inst_req_0); -- 
    cr_6338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2485_inst_req_1); -- 
    rr_6319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2481_inst_req_0); -- 
    cr_6324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2481_inst_req_1); -- 
    rr_6333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2485_inst_req_0); -- 
    cr_6310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2477_inst_req_1); -- 
    rr_6347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2515_inst_req_0); -- 
    cr_6352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2515_inst_req_1); -- 
    req_6383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => array_obj_ref_2521_index_offset_req_1); -- 
    req_6398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => addr_of_2522_final_reg_req_1); -- 
    cr_6443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => ptr_deref_2526_load_0_req_1); -- 
    req_6479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => array_obj_ref_2544_index_offset_req_1); -- 
    req_6494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => addr_of_2545_final_reg_req_1); -- 
    cr_6544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => ptr_deref_2548_store_0_req_1); -- 
    rr_6553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2553_inst_req_0); -- 
    cr_6558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(167), ack => type_cast_2553_inst_req_1); -- 
    convTransposeB_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(163) & convTransposeB_CP_5537_elements(164) & convTransposeB_CP_5537_elements(165) & convTransposeB_CP_5537_elements(166);
      gj_convTransposeB_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  transition  output  delay-element  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	139 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	175 
    -- CP-element group 168:  members (4) 
      -- CP-element group 168: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2628/$exit
      -- CP-element group 168: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/$exit
      -- CP-element group 168: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2632_konst_delay_trans
      -- CP-element group 168: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_req
      -- 
    phi_stmt_2628_req_6853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2628_req_6853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(168), ack => phi_stmt_2628_req_0); -- 
    -- Element group convTransposeB_CP_5537_elements(168) is a control-delay.
    cp_element_168_delay: control_delay_element  generic map(name => " 168_delay", delay_value => 1)  port map(req => convTransposeB_CP_5537_elements(139), ack => convTransposeB_CP_5537_elements(168), clk => clk, reset =>reset);
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	139 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/Sample/ra
      -- 
    ra_6870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2638_inst_ack_0, ack => convTransposeB_CP_5537_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	139 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (2) 
      -- CP-element group 170: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/Update/ca
      -- 
    ca_6875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2638_inst_ack_1, ack => convTransposeB_CP_5537_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	175 
    -- CP-element group 171:  members (5) 
      -- CP-element group 171: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/$exit
      -- CP-element group 171: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/$exit
      -- CP-element group 171: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/$exit
      -- CP-element group 171: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2638/SplitProtocol/$exit
      -- CP-element group 171: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_req
      -- 
    phi_stmt_2635_req_6876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2635_req_6876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(171), ack => phi_stmt_2635_req_0); -- 
    convTransposeB_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(169) & convTransposeB_CP_5537_elements(170);
      gj_convTransposeB_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	139 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/Sample/ra
      -- 
    ra_6893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2644_inst_ack_0, ack => convTransposeB_CP_5537_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	139 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (2) 
      -- CP-element group 173: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/Update/ca
      -- 
    ca_6898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2644_inst_ack_1, ack => convTransposeB_CP_5537_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/$exit
      -- CP-element group 174: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/$exit
      -- CP-element group 174: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/$exit
      -- CP-element group 174: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2644/SplitProtocol/$exit
      -- CP-element group 174: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_req
      -- 
    phi_stmt_2641_req_6899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2641_req_6899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(174), ack => phi_stmt_2641_req_0); -- 
    convTransposeB_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(172) & convTransposeB_CP_5537_elements(173);
      gj_convTransposeB_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: 	168 
    -- CP-element group 175: 	171 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	186 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_2070/ifx_xelse_ifx_xend254_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(174) & convTransposeB_CP_5537_elements(168) & convTransposeB_CP_5537_elements(171);
      gj_convTransposeB_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	130 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/Sample/ra
      -- 
    ra_6919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2634_inst_ack_0, ack => convTransposeB_CP_5537_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	130 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (2) 
      -- CP-element group 177: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/Update/ca
      -- 
    ca_6924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2634_inst_ack_1, ack => convTransposeB_CP_5537_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	185 
    -- CP-element group 178:  members (5) 
      -- CP-element group 178: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/$exit
      -- CP-element group 178: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/$exit
      -- CP-element group 178: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/$exit
      -- CP-element group 178: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_sources/type_cast_2634/SplitProtocol/$exit
      -- CP-element group 178: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2628/phi_stmt_2628_req
      -- 
    phi_stmt_2628_req_6925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2628_req_6925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(178), ack => phi_stmt_2628_req_1); -- 
    convTransposeB_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(176) & convTransposeB_CP_5537_elements(177);
      gj_convTransposeB_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	130 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/Sample/ra
      -- 
    ra_6942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2640_inst_ack_0, ack => convTransposeB_CP_5537_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	130 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/Update/ca
      -- 
    ca_6947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2640_inst_ack_1, ack => convTransposeB_CP_5537_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	185 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/$exit
      -- CP-element group 181: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/$exit
      -- CP-element group 181: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/$exit
      -- CP-element group 181: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_sources/type_cast_2640/SplitProtocol/$exit
      -- CP-element group 181: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2635/phi_stmt_2635_req
      -- 
    phi_stmt_2635_req_6948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2635_req_6948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(181), ack => phi_stmt_2635_req_1); -- 
    convTransposeB_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(179) & convTransposeB_CP_5537_elements(180);
      gj_convTransposeB_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	130 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/Sample/ra
      -- 
    ra_6965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2646_inst_ack_0, ack => convTransposeB_CP_5537_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	130 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/Update/ca
      -- 
    ca_6970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2646_inst_ack_1, ack => convTransposeB_CP_5537_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (5) 
      -- CP-element group 184: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/$exit
      -- CP-element group 184: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/$exit
      -- CP-element group 184: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/$exit
      -- CP-element group 184: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_sources/type_cast_2646/SplitProtocol/$exit
      -- CP-element group 184: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/phi_stmt_2641/phi_stmt_2641_req
      -- 
    phi_stmt_2641_req_6971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2641_req_6971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5537_elements(184), ack => phi_stmt_2641_req_1); -- 
    convTransposeB_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(182) & convTransposeB_CP_5537_elements(183);
      gj_convTransposeB_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	181 
    -- CP-element group 185: 	184 
    -- CP-element group 185: 	178 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_2070/ifx_xthen_ifx_xend254_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(181) & convTransposeB_CP_5537_elements(184) & convTransposeB_CP_5537_elements(178);
      gj_convTransposeB_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  merge  fork  transition  place  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	175 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	188 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (2) 
      -- CP-element group 186: 	 branch_block_stmt_2070/merge_stmt_2627_PhiReqMerge
      -- CP-element group 186: 	 branch_block_stmt_2070/merge_stmt_2627_PhiAck/$entry
      -- 
    convTransposeB_CP_5537_elements(186) <= OrReduce(convTransposeB_CP_5537_elements(175) & convTransposeB_CP_5537_elements(185));
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	190 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_2070/merge_stmt_2627_PhiAck/phi_stmt_2628_ack
      -- 
    phi_stmt_2628_ack_6976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2628_ack_0, ack => convTransposeB_CP_5537_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_2070/merge_stmt_2627_PhiAck/phi_stmt_2635_ack
      -- 
    phi_stmt_2635_ack_6977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2635_ack_0, ack => convTransposeB_CP_5537_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (1) 
      -- CP-element group 189: 	 branch_block_stmt_2070/merge_stmt_2627_PhiAck/phi_stmt_2641_ack
      -- 
    phi_stmt_2641_ack_6978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2641_ack_0, ack => convTransposeB_CP_5537_elements(189)); -- 
    -- CP-element group 190:  join  transition  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	187 
    -- CP-element group 190: 	188 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	1 
    -- CP-element group 190:  members (1) 
      -- CP-element group 190: 	 branch_block_stmt_2070/merge_stmt_2627_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_5537_elements(187) & convTransposeB_CP_5537_elements(188) & convTransposeB_CP_5537_elements(189);
      gj_convTransposeB_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5537_elements(190), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom212_2543_resized : std_logic_vector(13 downto 0);
    signal R_idxprom212_2543_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2520_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2520_scaled : std_logic_vector(13 downto 0);
    signal add103_2282 : std_logic_vector(31 downto 0);
    signal add108_2300 : std_logic_vector(31 downto 0);
    signal add113_2318 : std_logic_vector(31 downto 0);
    signal add135_2349 : std_logic_vector(63 downto 0);
    signal add147_2374 : std_logic_vector(63 downto 0);
    signal add16_2120 : std_logic_vector(31 downto 0);
    signal add171_2387 : std_logic_vector(15 downto 0);
    signal add184_2398 : std_logic_vector(15 downto 0);
    signal add203_2496 : std_logic_vector(63 downto 0);
    signal add205_2506 : std_logic_vector(63 downto 0);
    signal add217_2560 : std_logic_vector(31 downto 0);
    signal add224_2578 : std_logic_vector(15 downto 0);
    signal add28_2145 : std_logic_vector(31 downto 0);
    signal add52_2176 : std_logic_vector(15 downto 0);
    signal add64_2201 : std_logic_vector(15 downto 0);
    signal add86_2232 : std_logic_vector(15 downto 0);
    signal add95_2257 : std_logic_vector(15 downto 0);
    signal add_2095 : std_logic_vector(15 downto 0);
    signal add_src_0x_x0_2454 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2521_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2521_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2521_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2521_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2521_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2521_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2544_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2544_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2544_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2544_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2544_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2544_root_address : std_logic_vector(13 downto 0);
    signal arrayidx208_2523 : std_logic_vector(31 downto 0);
    signal arrayidx213_2546 : std_logic_vector(31 downto 0);
    signal call101_2273 : std_logic_vector(7 downto 0);
    signal call106_2291 : std_logic_vector(7 downto 0);
    signal call111_2309 : std_logic_vector(7 downto 0);
    signal call114_2321 : std_logic_vector(7 downto 0);
    signal call121_2324 : std_logic_vector(7 downto 0);
    signal call126_2327 : std_logic_vector(7 downto 0);
    signal call133_2340 : std_logic_vector(7 downto 0);
    signal call138_2352 : std_logic_vector(7 downto 0);
    signal call145_2365 : std_logic_vector(7 downto 0);
    signal call14_2111 : std_logic_vector(7 downto 0);
    signal call19_2123 : std_logic_vector(7 downto 0);
    signal call26_2136 : std_logic_vector(7 downto 0);
    signal call31_2148 : std_logic_vector(7 downto 0);
    signal call38_2151 : std_logic_vector(7 downto 0);
    signal call3_2086 : std_logic_vector(7 downto 0);
    signal call43_2154 : std_logic_vector(7 downto 0);
    signal call50_2167 : std_logic_vector(7 downto 0);
    signal call55_2179 : std_logic_vector(7 downto 0);
    signal call62_2192 : std_logic_vector(7 downto 0);
    signal call67_2204 : std_logic_vector(7 downto 0);
    signal call74_2207 : std_logic_vector(7 downto 0);
    signal call79_2210 : std_logic_vector(7 downto 0);
    signal call7_2098 : std_logic_vector(7 downto 0);
    signal call84_2223 : std_logic_vector(7 downto 0);
    signal call88_2235 : std_logic_vector(7 downto 0);
    signal call93_2248 : std_logic_vector(7 downto 0);
    signal call97_2260 : std_logic_vector(7 downto 0);
    signal call_2073 : std_logic_vector(7 downto 0);
    signal cmp232_2595 : std_logic_vector(0 downto 0);
    signal cmp243_2620 : std_logic_vector(0 downto 0);
    signal cmp_2565 : std_logic_vector(0 downto 0);
    signal conv102_2277 : std_logic_vector(31 downto 0);
    signal conv107_2295 : std_logic_vector(31 downto 0);
    signal conv112_2313 : std_logic_vector(31 downto 0);
    signal conv12_2102 : std_logic_vector(31 downto 0);
    signal conv131_2331 : std_logic_vector(63 downto 0);
    signal conv134_2344 : std_logic_vector(63 downto 0);
    signal conv143_2356 : std_logic_vector(63 downto 0);
    signal conv146_2369 : std_logic_vector(63 downto 0);
    signal conv15_2115 : std_logic_vector(31 downto 0);
    signal conv191_2478 : std_logic_vector(63 downto 0);
    signal conv196_2482 : std_logic_vector(63 downto 0);
    signal conv201_2486 : std_logic_vector(63 downto 0);
    signal conv216_2554 : std_logic_vector(31 downto 0);
    signal conv228_2590 : std_logic_vector(31 downto 0);
    signal conv238_2615 : std_logic_vector(31 downto 0);
    signal conv241_2407 : std_logic_vector(31 downto 0);
    signal conv24_2127 : std_logic_vector(31 downto 0);
    signal conv27_2140 : std_logic_vector(31 downto 0);
    signal conv2_2077 : std_logic_vector(15 downto 0);
    signal conv48_2158 : std_logic_vector(15 downto 0);
    signal conv4_2090 : std_logic_vector(15 downto 0);
    signal conv51_2171 : std_logic_vector(15 downto 0);
    signal conv60_2183 : std_logic_vector(15 downto 0);
    signal conv63_2196 : std_logic_vector(15 downto 0);
    signal conv82_2214 : std_logic_vector(15 downto 0);
    signal conv85_2227 : std_logic_vector(15 downto 0);
    signal conv91_2239 : std_logic_vector(15 downto 0);
    signal conv94_2252 : std_logic_vector(15 downto 0);
    signal conv98_2264 : std_logic_vector(31 downto 0);
    signal idxprom212_2539 : std_logic_vector(63 downto 0);
    signal idxprom_2516 : std_logic_vector(63 downto 0);
    signal inc236_2599 : std_logic_vector(15 downto 0);
    signal inc236x_xinput_dim0x_x2_2604 : std_logic_vector(15 downto 0);
    signal inc_2586 : std_logic_vector(15 downto 0);
    signal indvar_2416 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2653 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2641 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2437 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2635 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2430 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2611 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2628 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2423 : std_logic_vector(15 downto 0);
    signal mul180_2469 : std_logic_vector(15 downto 0);
    signal mul202_2491 : std_logic_vector(63 downto 0);
    signal mul204_2501 : std_logic_vector(63 downto 0);
    signal mul_2459 : std_logic_vector(15 downto 0);
    signal ptr_deref_2526_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2526_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2526_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2526_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2526_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2548_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2548_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2548_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2548_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2548_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2548_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl100_2270 : std_logic_vector(31 downto 0);
    signal shl105_2288 : std_logic_vector(31 downto 0);
    signal shl110_2306 : std_logic_vector(31 downto 0);
    signal shl132_2337 : std_logic_vector(63 downto 0);
    signal shl13_2108 : std_logic_vector(31 downto 0);
    signal shl144_2362 : std_logic_vector(63 downto 0);
    signal shl25_2133 : std_logic_vector(31 downto 0);
    signal shl49_2164 : std_logic_vector(15 downto 0);
    signal shl61_2189 : std_logic_vector(15 downto 0);
    signal shl83_2220 : std_logic_vector(15 downto 0);
    signal shl92_2245 : std_logic_vector(15 downto 0);
    signal shl_2083 : std_logic_vector(15 downto 0);
    signal shr207_2512 : std_logic_vector(31 downto 0);
    signal shr211_2533 : std_logic_vector(63 downto 0);
    signal shr242258_2413 : std_logic_vector(31 downto 0);
    signal shr257_2381 : std_logic_vector(15 downto 0);
    signal sub174_2464 : std_logic_vector(15 downto 0);
    signal sub187_2403 : std_logic_vector(15 downto 0);
    signal sub188_2474 : std_logic_vector(15 downto 0);
    signal sub_2392 : std_logic_vector(15 downto 0);
    signal tmp1_2449 : std_logic_vector(31 downto 0);
    signal tmp209_2527 : std_logic_vector(63 downto 0);
    signal type_cast_2081_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2106_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2131_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2162_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2187_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2218_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2243_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2268_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2286_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2304_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2335_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2360_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2379_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2385_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2396_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2411_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2420_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2422_wire : std_logic_vector(31 downto 0);
    signal type_cast_2426_wire : std_logic_vector(15 downto 0);
    signal type_cast_2429_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2433_wire : std_logic_vector(15 downto 0);
    signal type_cast_2436_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2440_wire : std_logic_vector(15 downto 0);
    signal type_cast_2442_wire : std_logic_vector(15 downto 0);
    signal type_cast_2447_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2510_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2531_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2537_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2558_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2576_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2584_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2608_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2632_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2634_wire : std_logic_vector(15 downto 0);
    signal type_cast_2638_wire : std_logic_vector(15 downto 0);
    signal type_cast_2640_wire : std_logic_vector(15 downto 0);
    signal type_cast_2644_wire : std_logic_vector(15 downto 0);
    signal type_cast_2646_wire : std_logic_vector(15 downto 0);
    signal type_cast_2651_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2659_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_2521_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2521_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2521_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2521_resized_base_address <= "00000000000000";
    array_obj_ref_2544_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2544_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2544_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2544_resized_base_address <= "00000000000000";
    ptr_deref_2526_word_offset_0 <= "00000000000000";
    ptr_deref_2548_word_offset_0 <= "00000000000000";
    type_cast_2081_wire_constant <= "0000000000001000";
    type_cast_2106_wire_constant <= "00000000000000000000000000001000";
    type_cast_2131_wire_constant <= "00000000000000000000000000001000";
    type_cast_2162_wire_constant <= "0000000000001000";
    type_cast_2187_wire_constant <= "0000000000001000";
    type_cast_2218_wire_constant <= "0000000000001000";
    type_cast_2243_wire_constant <= "0000000000001000";
    type_cast_2268_wire_constant <= "00000000000000000000000000001000";
    type_cast_2286_wire_constant <= "00000000000000000000000000001000";
    type_cast_2304_wire_constant <= "00000000000000000000000000001000";
    type_cast_2335_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2360_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2379_wire_constant <= "0000000000000010";
    type_cast_2385_wire_constant <= "1111111111111111";
    type_cast_2396_wire_constant <= "1111111111111111";
    type_cast_2411_wire_constant <= "00000000000000000000000000000001";
    type_cast_2420_wire_constant <= "00000000000000000000000000000000";
    type_cast_2429_wire_constant <= "0000000000000000";
    type_cast_2436_wire_constant <= "0000000000000000";
    type_cast_2447_wire_constant <= "00000000000000000000000000000100";
    type_cast_2510_wire_constant <= "00000000000000000000000000000010";
    type_cast_2531_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2537_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2558_wire_constant <= "00000000000000000000000000000100";
    type_cast_2576_wire_constant <= "0000000000000100";
    type_cast_2584_wire_constant <= "0000000000000001";
    type_cast_2608_wire_constant <= "0000000000000000";
    type_cast_2632_wire_constant <= "0000000000000000";
    type_cast_2651_wire_constant <= "00000000000000000000000000000001";
    type_cast_2659_wire_constant <= "00000001";
    phi_stmt_2416: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2420_wire_constant & type_cast_2422_wire;
      req <= phi_stmt_2416_req_0 & phi_stmt_2416_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2416",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2416_ack_0,
          idata => idata,
          odata => indvar_2416,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2416
    phi_stmt_2423: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2426_wire & type_cast_2429_wire_constant;
      req <= phi_stmt_2423_req_0 & phi_stmt_2423_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2423",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2423_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2423,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2423
    phi_stmt_2430: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2433_wire & type_cast_2436_wire_constant;
      req <= phi_stmt_2430_req_0 & phi_stmt_2430_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2430",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2430_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2430,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2430
    phi_stmt_2437: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2440_wire & type_cast_2442_wire;
      req <= phi_stmt_2437_req_0 & phi_stmt_2437_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2437",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2437_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2437,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2437
    phi_stmt_2628: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2632_wire_constant & type_cast_2634_wire;
      req <= phi_stmt_2628_req_0 & phi_stmt_2628_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2628",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2628_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2628,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2628
    phi_stmt_2635: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2638_wire & type_cast_2640_wire;
      req <= phi_stmt_2635_req_0 & phi_stmt_2635_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2635",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2635_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2635,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2635
    phi_stmt_2641: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2644_wire & type_cast_2646_wire;
      req <= phi_stmt_2641_req_0 & phi_stmt_2641_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2641",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2641_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2641,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2641
    -- flow-through select operator MUX_2610_inst
    input_dim1x_x2_2611 <= type_cast_2608_wire_constant when (cmp232_2595(0) /=  '0') else inc_2586;
    addr_of_2522_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2522_final_reg_req_0;
      addr_of_2522_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2522_final_reg_req_1;
      addr_of_2522_final_reg_ack_1<= rack(0);
      addr_of_2522_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2522_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2521_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx208_2523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2545_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2545_final_reg_req_0;
      addr_of_2545_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2545_final_reg_req_1;
      addr_of_2545_final_reg_ack_1<= rack(0);
      addr_of_2545_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2545_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2544_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx213_2546,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2076_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2076_inst_req_0;
      type_cast_2076_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2076_inst_req_1;
      type_cast_2076_inst_ack_1<= rack(0);
      type_cast_2076_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2076_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2073,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_2077,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2089_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2089_inst_req_0;
      type_cast_2089_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2089_inst_req_1;
      type_cast_2089_inst_ack_1<= rack(0);
      type_cast_2089_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2089_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2086,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_2090,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2101_inst_req_0;
      type_cast_2101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2101_inst_req_1;
      type_cast_2101_inst_ack_1<= rack(0);
      type_cast_2101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_2098,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_2102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2114_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2114_inst_req_0;
      type_cast_2114_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2114_inst_req_1;
      type_cast_2114_inst_ack_1<= rack(0);
      type_cast_2114_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2114_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_2111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_2115,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2126_inst_req_0;
      type_cast_2126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2126_inst_req_1;
      type_cast_2126_inst_ack_1<= rack(0);
      type_cast_2126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_2123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_2127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2139_inst_req_0;
      type_cast_2139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2139_inst_req_1;
      type_cast_2139_inst_ack_1<= rack(0);
      type_cast_2139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_2136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_2140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2157_inst_req_0;
      type_cast_2157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2157_inst_req_1;
      type_cast_2157_inst_ack_1<= rack(0);
      type_cast_2157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call43_2154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_2158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2170_inst_req_0;
      type_cast_2170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2170_inst_req_1;
      type_cast_2170_inst_ack_1<= rack(0);
      type_cast_2170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_2167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_2171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2182_inst_req_0;
      type_cast_2182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2182_inst_req_1;
      type_cast_2182_inst_ack_1<= rack(0);
      type_cast_2182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_2179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_2183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2195_inst_req_0;
      type_cast_2195_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2195_inst_req_1;
      type_cast_2195_inst_ack_1<= rack(0);
      type_cast_2195_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2195_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call62_2192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_2196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2213_inst_req_0;
      type_cast_2213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2213_inst_req_1;
      type_cast_2213_inst_ack_1<= rack(0);
      type_cast_2213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call79_2210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_2214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2226_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2226_inst_req_0;
      type_cast_2226_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2226_inst_req_1;
      type_cast_2226_inst_ack_1<= rack(0);
      type_cast_2226_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2226_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call84_2223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2227,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2238_inst_req_0;
      type_cast_2238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2238_inst_req_1;
      type_cast_2238_inst_ack_1<= rack(0);
      type_cast_2238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_2235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_2239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2251_inst_req_0;
      type_cast_2251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2251_inst_req_1;
      type_cast_2251_inst_ack_1<= rack(0);
      type_cast_2251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_2248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2263_inst_req_0;
      type_cast_2263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2263_inst_req_1;
      type_cast_2263_inst_ack_1<= rack(0);
      type_cast_2263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_2260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_2264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2276_inst_req_0;
      type_cast_2276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2276_inst_req_1;
      type_cast_2276_inst_ack_1<= rack(0);
      type_cast_2276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_2273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv102_2277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2294_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2294_inst_req_0;
      type_cast_2294_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2294_inst_req_1;
      type_cast_2294_inst_ack_1<= rack(0);
      type_cast_2294_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2294_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_2291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_2295,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2312_inst_req_0;
      type_cast_2312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2312_inst_req_1;
      type_cast_2312_inst_ack_1<= rack(0);
      type_cast_2312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_2309,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2330_inst_req_0;
      type_cast_2330_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2330_inst_req_1;
      type_cast_2330_inst_ack_1<= rack(0);
      type_cast_2330_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2330_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call126_2327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_2331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2343_inst_req_0;
      type_cast_2343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2343_inst_req_1;
      type_cast_2343_inst_ack_1<= rack(0);
      type_cast_2343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_2340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_2344,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2355_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2355_inst_req_0;
      type_cast_2355_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2355_inst_req_1;
      type_cast_2355_inst_ack_1<= rack(0);
      type_cast_2355_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2355_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call138_2352,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_2356,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2368_inst_req_0;
      type_cast_2368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2368_inst_req_1;
      type_cast_2368_inst_ack_1<= rack(0);
      type_cast_2368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_2365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv146_2369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2406_inst_req_0;
      type_cast_2406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2406_inst_req_1;
      type_cast_2406_inst_ack_1<= rack(0);
      type_cast_2406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_2095,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_2407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2422_inst_req_0;
      type_cast_2422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2422_inst_req_1;
      type_cast_2422_inst_ack_1<= rack(0);
      type_cast_2422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2422_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2426_inst_req_0;
      type_cast_2426_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2426_inst_req_1;
      type_cast_2426_inst_ack_1<= rack(0);
      type_cast_2426_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2426_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2426_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2433_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2433_inst_req_0;
      type_cast_2433_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2433_inst_req_1;
      type_cast_2433_inst_ack_1<= rack(0);
      type_cast_2433_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2433_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2635,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2433_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2440_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2440_inst_req_0;
      type_cast_2440_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2440_inst_req_1;
      type_cast_2440_inst_ack_1<= rack(0);
      type_cast_2440_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2440_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2440_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2442_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2442_inst_req_0;
      type_cast_2442_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2442_inst_req_1;
      type_cast_2442_inst_ack_1<= rack(0);
      type_cast_2442_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2442_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr257_2381,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2442_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2477_inst_req_0;
      type_cast_2477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2477_inst_req_1;
      type_cast_2477_inst_ack_1<= rack(0);
      type_cast_2477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_2478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2481_inst_req_0;
      type_cast_2481_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2481_inst_req_1;
      type_cast_2481_inst_ack_1<= rack(0);
      type_cast_2481_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2481_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub188_2474,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv196_2482,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2485_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2485_inst_req_0;
      type_cast_2485_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2485_inst_req_1;
      type_cast_2485_inst_ack_1<= rack(0);
      type_cast_2485_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2485_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub174_2464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv201_2486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2515_inst_req_0;
      type_cast_2515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2515_inst_req_1;
      type_cast_2515_inst_ack_1<= rack(0);
      type_cast_2515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr207_2512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2553_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2553_inst_req_0;
      type_cast_2553_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2553_inst_req_1;
      type_cast_2553_inst_ack_1<= rack(0);
      type_cast_2553_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2553_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv216_2554,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2589_inst_req_0;
      type_cast_2589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2589_inst_req_1;
      type_cast_2589_inst_ack_1<= rack(0);
      type_cast_2589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv228_2590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2598_inst_req_0;
      type_cast_2598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2598_inst_req_1;
      type_cast_2598_inst_ack_1<= rack(0);
      type_cast_2598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp232_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc236_2599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2614_inst_req_0;
      type_cast_2614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2614_inst_req_1;
      type_cast_2614_inst_ack_1<= rack(0);
      type_cast_2614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc236x_xinput_dim0x_x2_2604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv238_2615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2634_inst_req_0;
      type_cast_2634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2634_inst_req_1;
      type_cast_2634_inst_ack_1<= rack(0);
      type_cast_2634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add224_2578,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2634_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2638_inst_req_0;
      type_cast_2638_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2638_inst_req_1;
      type_cast_2638_inst_ack_1<= rack(0);
      type_cast_2638_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2638_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2638_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2640_inst_req_0;
      type_cast_2640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2640_inst_req_1;
      type_cast_2640_inst_ack_1<= rack(0);
      type_cast_2640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2430,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2640_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2644_inst_req_0;
      type_cast_2644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2644_inst_req_1;
      type_cast_2644_inst_ack_1<= rack(0);
      type_cast_2644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc236x_xinput_dim0x_x2_2604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2644_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2646_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2646_inst_req_0;
      type_cast_2646_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2646_inst_req_1;
      type_cast_2646_inst_ack_1<= rack(0);
      type_cast_2646_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2646_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2437,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2646_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2521_index_1_rename
    process(R_idxprom_2520_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2520_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2520_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2521_index_1_resize
    process(idxprom_2516) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2516;
      ov := iv(13 downto 0);
      R_idxprom_2520_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2521_root_address_inst
    process(array_obj_ref_2521_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2521_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2521_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2544_index_1_rename
    process(R_idxprom212_2543_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom212_2543_resized;
      ov(13 downto 0) := iv;
      R_idxprom212_2543_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2544_index_1_resize
    process(idxprom212_2539) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom212_2539;
      ov := iv(13 downto 0);
      R_idxprom212_2543_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2544_root_address_inst
    process(array_obj_ref_2544_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2544_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2544_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2526_addr_0
    process(ptr_deref_2526_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2526_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2526_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2526_base_resize
    process(arrayidx208_2523) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx208_2523;
      ov := iv(13 downto 0);
      ptr_deref_2526_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2526_gather_scatter
    process(ptr_deref_2526_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2526_data_0;
      ov(63 downto 0) := iv;
      tmp209_2527 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2526_root_address_inst
    process(ptr_deref_2526_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2526_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2526_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2548_addr_0
    process(ptr_deref_2548_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2548_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2548_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2548_base_resize
    process(arrayidx213_2546) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx213_2546;
      ov := iv(13 downto 0);
      ptr_deref_2548_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2548_gather_scatter
    process(tmp209_2527) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp209_2527;
      ov(63 downto 0) := iv;
      ptr_deref_2548_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2548_root_address_inst
    process(ptr_deref_2548_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2548_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2548_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2566_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2565;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2566_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2566_branch_req_0,
          ack0 => if_stmt_2566_branch_ack_0,
          ack1 => if_stmt_2566_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2621_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp243_2620;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2621_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2621_branch_req_0,
          ack0 => if_stmt_2621_branch_ack_0,
          ack1 => if_stmt_2621_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2386_inst
    process(add52_2176) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add52_2176, type_cast_2385_wire_constant, tmp_var);
      add171_2387 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2397_inst
    process(add64_2201) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add64_2201, type_cast_2396_wire_constant, tmp_var);
      add184_2398 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2463_inst
    process(sub_2392, mul_2459) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2392, mul_2459, tmp_var);
      sub174_2464 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2473_inst
    process(sub187_2403, mul180_2469) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub187_2403, mul180_2469, tmp_var);
      sub188_2474 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2577_inst
    process(input_dim2x_x1_2423) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2423, type_cast_2576_wire_constant, tmp_var);
      add224_2578 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2585_inst
    process(input_dim1x_x1_2430) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2430, type_cast_2584_wire_constant, tmp_var);
      inc_2586 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2603_inst
    process(inc236_2599, input_dim0x_x2_2437) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc236_2599, input_dim0x_x2_2437, tmp_var);
      inc236x_xinput_dim0x_x2_2604 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2453_inst
    process(add113_2318, tmp1_2449) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add113_2318, tmp1_2449, tmp_var);
      add_src_0x_x0_2454 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2559_inst
    process(conv216_2554) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv216_2554, type_cast_2558_wire_constant, tmp_var);
      add217_2560 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2652_inst
    process(indvar_2416) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2416, type_cast_2651_wire_constant, tmp_var);
      indvarx_xnext_2653 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2495_inst
    process(mul202_2491, conv196_2482) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul202_2491, conv196_2482, tmp_var);
      add203_2496 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2505_inst
    process(mul204_2501, conv191_2478) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul204_2501, conv191_2478, tmp_var);
      add205_2506 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2538_inst
    process(shr211_2533) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr211_2533, type_cast_2537_wire_constant, tmp_var);
      idxprom212_2539 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2594_inst
    process(conv228_2590, add16_2120) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv228_2590, add16_2120, tmp_var);
      cmp232_2595 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2619_inst
    process(conv238_2615, shr242258_2413) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv238_2615, shr242258_2413, tmp_var);
      cmp243_2620 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2380_inst
    process(add_2095) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_2095, type_cast_2379_wire_constant, tmp_var);
      shr257_2381 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2412_inst
    process(conv241_2407) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv241_2407, type_cast_2411_wire_constant, tmp_var);
      shr242258_2413 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2511_inst
    process(add_src_0x_x0_2454) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2454, type_cast_2510_wire_constant, tmp_var);
      shr207_2512 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2532_inst
    process(add205_2506) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add205_2506, type_cast_2531_wire_constant, tmp_var);
      shr211_2533 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2458_inst
    process(input_dim0x_x2_2437, add86_2232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2437, add86_2232, tmp_var);
      mul_2459 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2468_inst
    process(input_dim1x_x1_2430, add86_2232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2430, add86_2232, tmp_var);
      mul180_2469 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2448_inst
    process(indvar_2416) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2416, type_cast_2447_wire_constant, tmp_var);
      tmp1_2449 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2490_inst
    process(conv201_2486, add135_2349) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv201_2486, add135_2349, tmp_var);
      mul202_2491 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2500_inst
    process(add203_2496, add147_2374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add203_2496, add147_2374, tmp_var);
      mul204_2501 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2094_inst
    process(shl_2083, conv4_2090) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2083, conv4_2090, tmp_var);
      add_2095 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2175_inst
    process(shl49_2164, conv51_2171) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl49_2164, conv51_2171, tmp_var);
      add52_2176 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2200_inst
    process(shl61_2189, conv63_2196) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl61_2189, conv63_2196, tmp_var);
      add64_2201 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2231_inst
    process(shl83_2220, conv85_2227) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl83_2220, conv85_2227, tmp_var);
      add86_2232 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2256_inst
    process(shl92_2245, conv94_2252) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_2245, conv94_2252, tmp_var);
      add95_2257 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2119_inst
    process(shl13_2108, conv15_2115) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl13_2108, conv15_2115, tmp_var);
      add16_2120 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2144_inst
    process(shl25_2133, conv27_2140) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl25_2133, conv27_2140, tmp_var);
      add28_2145 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2281_inst
    process(shl100_2270, conv102_2277) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_2270, conv102_2277, tmp_var);
      add103_2282 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2299_inst
    process(shl105_2288, conv107_2295) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_2288, conv107_2295, tmp_var);
      add108_2300 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2317_inst
    process(shl110_2306, conv112_2313) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_2306, conv112_2313, tmp_var);
      add113_2318 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2348_inst
    process(shl132_2337, conv134_2344) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_2337, conv134_2344, tmp_var);
      add135_2349 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2373_inst
    process(shl144_2362, conv146_2369) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_2362, conv146_2369, tmp_var);
      add147_2374 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2082_inst
    process(conv2_2077) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv2_2077, type_cast_2081_wire_constant, tmp_var);
      shl_2083 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2163_inst
    process(conv48_2158) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_2158, type_cast_2162_wire_constant, tmp_var);
      shl49_2164 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2188_inst
    process(conv60_2183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv60_2183, type_cast_2187_wire_constant, tmp_var);
      shl61_2189 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2219_inst
    process(conv82_2214) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv82_2214, type_cast_2218_wire_constant, tmp_var);
      shl83_2220 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2244_inst
    process(conv91_2239) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_2239, type_cast_2243_wire_constant, tmp_var);
      shl92_2245 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2107_inst
    process(conv12_2102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv12_2102, type_cast_2106_wire_constant, tmp_var);
      shl13_2108 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2132_inst
    process(conv24_2127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv24_2127, type_cast_2131_wire_constant, tmp_var);
      shl25_2133 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2269_inst
    process(conv98_2264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv98_2264, type_cast_2268_wire_constant, tmp_var);
      shl100_2270 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2287_inst
    process(add103_2282) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add103_2282, type_cast_2286_wire_constant, tmp_var);
      shl105_2288 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2305_inst
    process(add108_2300) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_2300, type_cast_2304_wire_constant, tmp_var);
      shl110_2306 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2336_inst
    process(conv131_2331) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_2331, type_cast_2335_wire_constant, tmp_var);
      shl132_2337 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2361_inst
    process(conv143_2356) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv143_2356, type_cast_2360_wire_constant, tmp_var);
      shl144_2362 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2391_inst
    process(add171_2387, add95_2257) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add171_2387, add95_2257, tmp_var);
      sub_2392 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2402_inst
    process(add184_2398, add95_2257) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add184_2398, add95_2257, tmp_var);
      sub187_2403 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2564_inst
    process(add217_2560, add28_2145) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add217_2560, add28_2145, tmp_var);
      cmp_2565 <= tmp_var; --
    end process;
    -- shared split operator group (51) : array_obj_ref_2521_index_offset 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2520_scaled;
      array_obj_ref_2521_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2521_index_offset_req_0;
      array_obj_ref_2521_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2521_index_offset_req_1;
      array_obj_ref_2521_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : array_obj_ref_2544_index_offset 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom212_2543_scaled;
      array_obj_ref_2544_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2544_index_offset_req_0;
      array_obj_ref_2544_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2544_index_offset_req_1;
      array_obj_ref_2544_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared load operator group (0) : ptr_deref_2526_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2526_load_0_req_0;
      ptr_deref_2526_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2526_load_0_req_1;
      ptr_deref_2526_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2526_word_address_0;
      ptr_deref_2526_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2548_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2548_store_0_req_0;
      ptr_deref_2548_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2548_store_0_req_1;
      ptr_deref_2548_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2548_word_address_0;
      data_in <= ptr_deref_2548_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_2135_inst RPIPE_Block1_start_2272_inst RPIPE_Block1_start_2364_inst RPIPE_Block1_start_2147_inst RPIPE_Block1_start_2339_inst RPIPE_Block1_start_2150_inst RPIPE_Block1_start_2153_inst RPIPE_Block1_start_2166_inst RPIPE_Block1_start_2326_inst RPIPE_Block1_start_2351_inst RPIPE_Block1_start_2323_inst RPIPE_Block1_start_2320_inst RPIPE_Block1_start_2122_inst RPIPE_Block1_start_2247_inst RPIPE_Block1_start_2290_inst RPIPE_Block1_start_2259_inst RPIPE_Block1_start_2110_inst RPIPE_Block1_start_2234_inst RPIPE_Block1_start_2222_inst RPIPE_Block1_start_2097_inst RPIPE_Block1_start_2209_inst RPIPE_Block1_start_2085_inst RPIPE_Block1_start_2206_inst RPIPE_Block1_start_2308_inst RPIPE_Block1_start_2203_inst RPIPE_Block1_start_2191_inst RPIPE_Block1_start_2178_inst RPIPE_Block1_start_2072_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 27 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 27 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant outBUFs : IntegerArray(27 downto 0) := (27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      reqL_unguarded(27) <= RPIPE_Block1_start_2135_inst_req_0;
      reqL_unguarded(26) <= RPIPE_Block1_start_2272_inst_req_0;
      reqL_unguarded(25) <= RPIPE_Block1_start_2364_inst_req_0;
      reqL_unguarded(24) <= RPIPE_Block1_start_2147_inst_req_0;
      reqL_unguarded(23) <= RPIPE_Block1_start_2339_inst_req_0;
      reqL_unguarded(22) <= RPIPE_Block1_start_2150_inst_req_0;
      reqL_unguarded(21) <= RPIPE_Block1_start_2153_inst_req_0;
      reqL_unguarded(20) <= RPIPE_Block1_start_2166_inst_req_0;
      reqL_unguarded(19) <= RPIPE_Block1_start_2326_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Block1_start_2351_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Block1_start_2323_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Block1_start_2320_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Block1_start_2122_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Block1_start_2247_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Block1_start_2290_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_2259_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_2110_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_2234_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_2222_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_2097_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_2209_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_2085_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_2206_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_2308_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_2203_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_2191_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_2178_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_2072_inst_req_0;
      RPIPE_Block1_start_2135_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_Block1_start_2272_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_Block1_start_2364_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_Block1_start_2147_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_Block1_start_2339_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_Block1_start_2150_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_Block1_start_2153_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_Block1_start_2166_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_Block1_start_2326_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Block1_start_2351_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Block1_start_2323_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Block1_start_2320_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Block1_start_2122_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Block1_start_2247_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Block1_start_2290_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_2259_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_2110_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_2234_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_2222_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_2097_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_2209_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_2085_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_2206_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_2308_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_2203_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_2191_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_2178_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_2072_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(27) <= RPIPE_Block1_start_2135_inst_req_1;
      reqR_unguarded(26) <= RPIPE_Block1_start_2272_inst_req_1;
      reqR_unguarded(25) <= RPIPE_Block1_start_2364_inst_req_1;
      reqR_unguarded(24) <= RPIPE_Block1_start_2147_inst_req_1;
      reqR_unguarded(23) <= RPIPE_Block1_start_2339_inst_req_1;
      reqR_unguarded(22) <= RPIPE_Block1_start_2150_inst_req_1;
      reqR_unguarded(21) <= RPIPE_Block1_start_2153_inst_req_1;
      reqR_unguarded(20) <= RPIPE_Block1_start_2166_inst_req_1;
      reqR_unguarded(19) <= RPIPE_Block1_start_2326_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Block1_start_2351_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Block1_start_2323_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Block1_start_2320_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Block1_start_2122_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Block1_start_2247_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Block1_start_2290_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_2259_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_2110_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_2234_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_2222_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_2097_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_2209_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_2085_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_2206_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_2308_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_2203_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_2191_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_2178_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_2072_inst_req_1;
      RPIPE_Block1_start_2135_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_Block1_start_2272_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_Block1_start_2364_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_Block1_start_2147_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_Block1_start_2339_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_Block1_start_2150_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_Block1_start_2153_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_Block1_start_2166_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_Block1_start_2326_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Block1_start_2351_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Block1_start_2323_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Block1_start_2320_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Block1_start_2122_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Block1_start_2247_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Block1_start_2290_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_2259_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_2110_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_2234_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_2222_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_2097_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_2209_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_2085_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_2206_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_2308_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_2203_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_2191_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_2178_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_2072_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      call26_2136 <= data_out(223 downto 216);
      call101_2273 <= data_out(215 downto 208);
      call145_2365 <= data_out(207 downto 200);
      call31_2148 <= data_out(199 downto 192);
      call133_2340 <= data_out(191 downto 184);
      call38_2151 <= data_out(183 downto 176);
      call43_2154 <= data_out(175 downto 168);
      call50_2167 <= data_out(167 downto 160);
      call126_2327 <= data_out(159 downto 152);
      call138_2352 <= data_out(151 downto 144);
      call121_2324 <= data_out(143 downto 136);
      call114_2321 <= data_out(135 downto 128);
      call19_2123 <= data_out(127 downto 120);
      call93_2248 <= data_out(119 downto 112);
      call106_2291 <= data_out(111 downto 104);
      call97_2260 <= data_out(103 downto 96);
      call14_2111 <= data_out(95 downto 88);
      call88_2235 <= data_out(87 downto 80);
      call84_2223 <= data_out(79 downto 72);
      call7_2098 <= data_out(71 downto 64);
      call79_2210 <= data_out(63 downto 56);
      call3_2086 <= data_out(55 downto 48);
      call74_2207 <= data_out(47 downto 40);
      call111_2309 <= data_out(39 downto 32);
      call67_2204 <= data_out(31 downto 24);
      call62_2192 <= data_out(23 downto 16);
      call55_2179 <= data_out(15 downto 8);
      call_2073 <= data_out(7 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 8,  num_reqs => 28,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2657_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2657_inst_req_0;
      WPIPE_Block1_done_2657_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2657_inst_req_1;
      WPIPE_Block1_done_2657_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2659_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_6995_start: Boolean;
  signal convTransposeC_CP_6995_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_3092_inst_ack_0 : boolean;
  signal type_cast_3084_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2947_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2947_inst_ack_0 : boolean;
  signal type_cast_2951_inst_req_0 : boolean;
  signal type_cast_3092_inst_req_0 : boolean;
  signal type_cast_2964_inst_req_1 : boolean;
  signal type_cast_2926_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2947_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2935_inst_ack_0 : boolean;
  signal type_cast_2951_inst_ack_0 : boolean;
  signal type_cast_2926_inst_ack_0 : boolean;
  signal type_cast_2964_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2960_inst_req_1 : boolean;
  signal type_cast_3002_inst_req_0 : boolean;
  signal type_cast_3122_inst_req_0 : boolean;
  signal type_cast_3084_inst_req_0 : boolean;
  signal type_cast_3002_inst_ack_0 : boolean;
  signal type_cast_2964_inst_req_0 : boolean;
  signal array_obj_ref_3128_index_offset_ack_0 : boolean;
  signal type_cast_2964_inst_ack_1 : boolean;
  signal type_cast_3088_inst_ack_1 : boolean;
  signal type_cast_3088_inst_req_1 : boolean;
  signal type_cast_3122_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2935_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2935_inst_req_1 : boolean;
  signal type_cast_2939_inst_req_0 : boolean;
  signal type_cast_2926_inst_req_0 : boolean;
  signal type_cast_3122_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2960_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2947_inst_ack_1 : boolean;
  signal type_cast_3122_inst_ack_0 : boolean;
  signal type_cast_2939_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2935_inst_req_0 : boolean;
  signal type_cast_3088_inst_ack_0 : boolean;
  signal array_obj_ref_3128_index_offset_ack_1 : boolean;
  signal type_cast_3088_inst_req_0 : boolean;
  signal addr_of_3129_final_reg_ack_1 : boolean;
  signal RPIPE_Block2_start_2922_inst_ack_1 : boolean;
  signal type_cast_2926_inst_ack_1 : boolean;
  signal array_obj_ref_3128_index_offset_req_1 : boolean;
  signal type_cast_2951_inst_req_1 : boolean;
  signal ptr_deref_3133_load_0_ack_1 : boolean;
  signal addr_of_3152_final_reg_req_1 : boolean;
  signal ptr_deref_3133_load_0_ack_0 : boolean;
  signal type_cast_2951_inst_ack_1 : boolean;
  signal type_cast_3002_inst_req_1 : boolean;
  signal addr_of_3152_final_reg_req_0 : boolean;
  signal type_cast_2939_inst_ack_0 : boolean;
  signal addr_of_3129_final_reg_req_0 : boolean;
  signal array_obj_ref_3151_index_offset_req_1 : boolean;
  signal addr_of_3152_final_reg_ack_0 : boolean;
  signal addr_of_3129_final_reg_ack_0 : boolean;
  signal type_cast_3002_inst_ack_1 : boolean;
  signal type_cast_3092_inst_req_1 : boolean;
  signal type_cast_3092_inst_ack_1 : boolean;
  signal type_cast_3084_inst_req_1 : boolean;
  signal type_cast_3084_inst_ack_1 : boolean;
  signal array_obj_ref_3151_index_offset_req_0 : boolean;
  signal type_cast_2939_inst_req_1 : boolean;
  signal array_obj_ref_3151_index_offset_ack_1 : boolean;
  signal ptr_deref_3133_load_0_req_1 : boolean;
  signal RPIPE_Block2_start_2960_inst_req_0 : boolean;
  signal array_obj_ref_3151_index_offset_ack_0 : boolean;
  signal RPIPE_Block2_start_2960_inst_ack_0 : boolean;
  signal array_obj_ref_3128_index_offset_req_0 : boolean;
  signal addr_of_3129_final_reg_req_1 : boolean;
  signal ptr_deref_3133_load_0_req_0 : boolean;
  signal RPIPE_Block2_start_2922_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2668_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2668_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2668_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2668_inst_ack_1 : boolean;
  signal type_cast_2672_inst_req_0 : boolean;
  signal type_cast_2672_inst_ack_0 : boolean;
  signal type_cast_2672_inst_req_1 : boolean;
  signal type_cast_2672_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2681_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2681_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2681_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2681_inst_ack_1 : boolean;
  signal type_cast_2685_inst_req_0 : boolean;
  signal type_cast_2685_inst_ack_0 : boolean;
  signal type_cast_2685_inst_req_1 : boolean;
  signal type_cast_2685_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2693_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2693_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2693_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2693_inst_ack_1 : boolean;
  signal type_cast_2697_inst_req_0 : boolean;
  signal type_cast_2697_inst_ack_0 : boolean;
  signal type_cast_2697_inst_req_1 : boolean;
  signal type_cast_2697_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2706_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2706_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2706_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2706_inst_ack_1 : boolean;
  signal type_cast_2710_inst_req_0 : boolean;
  signal type_cast_2710_inst_ack_0 : boolean;
  signal type_cast_2710_inst_req_1 : boolean;
  signal type_cast_2710_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2718_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2718_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2718_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2718_inst_ack_1 : boolean;
  signal type_cast_2722_inst_req_0 : boolean;
  signal type_cast_2722_inst_ack_0 : boolean;
  signal type_cast_2722_inst_req_1 : boolean;
  signal type_cast_2722_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2731_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2731_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2731_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2731_inst_ack_1 : boolean;
  signal type_cast_2735_inst_req_0 : boolean;
  signal type_cast_2735_inst_ack_0 : boolean;
  signal type_cast_2735_inst_req_1 : boolean;
  signal type_cast_2735_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2743_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2743_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2743_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2743_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2746_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2746_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2746_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2746_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2749_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2749_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2749_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2749_inst_ack_1 : boolean;
  signal type_cast_2753_inst_req_0 : boolean;
  signal type_cast_2753_inst_ack_0 : boolean;
  signal type_cast_2753_inst_req_1 : boolean;
  signal type_cast_2753_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2762_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2762_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2762_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2762_inst_ack_1 : boolean;
  signal type_cast_2766_inst_req_0 : boolean;
  signal type_cast_2766_inst_ack_0 : boolean;
  signal type_cast_2766_inst_req_1 : boolean;
  signal type_cast_2766_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2774_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2774_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2774_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2774_inst_ack_1 : boolean;
  signal type_cast_2778_inst_req_0 : boolean;
  signal type_cast_2778_inst_ack_0 : boolean;
  signal type_cast_2778_inst_req_1 : boolean;
  signal type_cast_2778_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2787_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2787_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2787_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2787_inst_ack_1 : boolean;
  signal addr_of_3152_final_reg_ack_1 : boolean;
  signal type_cast_2791_inst_req_0 : boolean;
  signal type_cast_2791_inst_ack_0 : boolean;
  signal type_cast_2791_inst_req_1 : boolean;
  signal type_cast_2791_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2799_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2799_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2799_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2799_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2802_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2802_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2802_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2802_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2805_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2805_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2805_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2805_inst_ack_1 : boolean;
  signal type_cast_2809_inst_req_0 : boolean;
  signal type_cast_2809_inst_ack_0 : boolean;
  signal type_cast_2809_inst_req_1 : boolean;
  signal type_cast_2809_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2818_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2818_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2818_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2818_inst_ack_1 : boolean;
  signal type_cast_2822_inst_req_0 : boolean;
  signal type_cast_2822_inst_ack_0 : boolean;
  signal type_cast_2822_inst_req_1 : boolean;
  signal type_cast_2822_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2830_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2830_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2830_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2830_inst_ack_1 : boolean;
  signal type_cast_2834_inst_req_0 : boolean;
  signal type_cast_2834_inst_ack_0 : boolean;
  signal type_cast_2834_inst_req_1 : boolean;
  signal type_cast_2834_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2843_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2843_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2843_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2843_inst_ack_1 : boolean;
  signal type_cast_2847_inst_req_0 : boolean;
  signal type_cast_2847_inst_ack_0 : boolean;
  signal type_cast_2847_inst_req_1 : boolean;
  signal type_cast_2847_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2855_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2855_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2855_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2855_inst_ack_1 : boolean;
  signal type_cast_2859_inst_req_0 : boolean;
  signal type_cast_2859_inst_ack_0 : boolean;
  signal type_cast_2859_inst_req_1 : boolean;
  signal type_cast_2859_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2868_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2868_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2868_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2868_inst_ack_1 : boolean;
  signal type_cast_2872_inst_req_0 : boolean;
  signal type_cast_2872_inst_ack_0 : boolean;
  signal type_cast_2872_inst_req_1 : boolean;
  signal type_cast_2872_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2886_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2886_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2886_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2886_inst_ack_1 : boolean;
  signal type_cast_2890_inst_req_0 : boolean;
  signal type_cast_2890_inst_ack_0 : boolean;
  signal type_cast_2890_inst_req_1 : boolean;
  signal type_cast_2890_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2904_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2904_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2904_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2904_inst_ack_1 : boolean;
  signal type_cast_2908_inst_req_0 : boolean;
  signal type_cast_2908_inst_ack_0 : boolean;
  signal type_cast_2908_inst_req_1 : boolean;
  signal type_cast_2908_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2916_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2916_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2916_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2916_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2919_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2919_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2919_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2919_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2922_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2922_inst_ack_0 : boolean;
  signal ptr_deref_3155_store_0_req_0 : boolean;
  signal ptr_deref_3155_store_0_ack_0 : boolean;
  signal ptr_deref_3155_store_0_req_1 : boolean;
  signal ptr_deref_3155_store_0_ack_1 : boolean;
  signal type_cast_3160_inst_req_0 : boolean;
  signal type_cast_3160_inst_ack_0 : boolean;
  signal type_cast_3160_inst_req_1 : boolean;
  signal type_cast_3160_inst_ack_1 : boolean;
  signal if_stmt_3173_branch_req_0 : boolean;
  signal if_stmt_3173_branch_ack_1 : boolean;
  signal if_stmt_3173_branch_ack_0 : boolean;
  signal type_cast_3196_inst_req_0 : boolean;
  signal type_cast_3196_inst_ack_0 : boolean;
  signal type_cast_3196_inst_req_1 : boolean;
  signal type_cast_3196_inst_ack_1 : boolean;
  signal type_cast_3205_inst_req_0 : boolean;
  signal type_cast_3205_inst_ack_0 : boolean;
  signal type_cast_3205_inst_req_1 : boolean;
  signal type_cast_3205_inst_ack_1 : boolean;
  signal type_cast_3221_inst_req_0 : boolean;
  signal type_cast_3221_inst_ack_0 : boolean;
  signal type_cast_3221_inst_req_1 : boolean;
  signal type_cast_3221_inst_ack_1 : boolean;
  signal if_stmt_3228_branch_req_0 : boolean;
  signal if_stmt_3228_branch_ack_1 : boolean;
  signal if_stmt_3228_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_3264_inst_req_0 : boolean;
  signal WPIPE_Block2_done_3264_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_3264_inst_req_1 : boolean;
  signal WPIPE_Block2_done_3264_inst_ack_1 : boolean;
  signal phi_stmt_3023_req_0 : boolean;
  signal phi_stmt_3030_req_0 : boolean;
  signal phi_stmt_3037_req_0 : boolean;
  signal type_cast_3047_inst_req_0 : boolean;
  signal type_cast_3047_inst_ack_0 : boolean;
  signal type_cast_3047_inst_req_1 : boolean;
  signal type_cast_3047_inst_ack_1 : boolean;
  signal phi_stmt_3044_req_0 : boolean;
  signal type_cast_3029_inst_req_0 : boolean;
  signal type_cast_3029_inst_ack_0 : boolean;
  signal type_cast_3029_inst_req_1 : boolean;
  signal type_cast_3029_inst_ack_1 : boolean;
  signal phi_stmt_3023_req_1 : boolean;
  signal type_cast_3036_inst_req_0 : boolean;
  signal type_cast_3036_inst_ack_0 : boolean;
  signal type_cast_3036_inst_req_1 : boolean;
  signal type_cast_3036_inst_ack_1 : boolean;
  signal phi_stmt_3030_req_1 : boolean;
  signal type_cast_3043_inst_req_0 : boolean;
  signal type_cast_3043_inst_ack_0 : boolean;
  signal type_cast_3043_inst_req_1 : boolean;
  signal type_cast_3043_inst_ack_1 : boolean;
  signal phi_stmt_3037_req_1 : boolean;
  signal type_cast_3049_inst_req_0 : boolean;
  signal type_cast_3049_inst_ack_0 : boolean;
  signal type_cast_3049_inst_req_1 : boolean;
  signal type_cast_3049_inst_ack_1 : boolean;
  signal phi_stmt_3044_req_1 : boolean;
  signal phi_stmt_3023_ack_0 : boolean;
  signal phi_stmt_3030_ack_0 : boolean;
  signal phi_stmt_3037_ack_0 : boolean;
  signal phi_stmt_3044_ack_0 : boolean;
  signal phi_stmt_3235_req_1 : boolean;
  signal type_cast_3247_inst_req_0 : boolean;
  signal type_cast_3247_inst_ack_0 : boolean;
  signal type_cast_3247_inst_req_1 : boolean;
  signal type_cast_3247_inst_ack_1 : boolean;
  signal phi_stmt_3242_req_1 : boolean;
  signal type_cast_3253_inst_req_0 : boolean;
  signal type_cast_3253_inst_ack_0 : boolean;
  signal type_cast_3253_inst_req_1 : boolean;
  signal type_cast_3253_inst_ack_1 : boolean;
  signal phi_stmt_3248_req_1 : boolean;
  signal type_cast_3238_inst_req_0 : boolean;
  signal type_cast_3238_inst_ack_0 : boolean;
  signal type_cast_3238_inst_req_1 : boolean;
  signal type_cast_3238_inst_ack_1 : boolean;
  signal phi_stmt_3235_req_0 : boolean;
  signal type_cast_3245_inst_req_0 : boolean;
  signal type_cast_3245_inst_ack_0 : boolean;
  signal type_cast_3245_inst_req_1 : boolean;
  signal type_cast_3245_inst_ack_1 : boolean;
  signal phi_stmt_3242_req_0 : boolean;
  signal type_cast_3251_inst_req_0 : boolean;
  signal type_cast_3251_inst_ack_0 : boolean;
  signal type_cast_3251_inst_req_1 : boolean;
  signal type_cast_3251_inst_ack_1 : boolean;
  signal phi_stmt_3248_req_0 : boolean;
  signal phi_stmt_3235_ack_0 : boolean;
  signal phi_stmt_3242_ack_0 : boolean;
  signal phi_stmt_3248_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_6995_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6995_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_6995_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6995_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_6995: Block -- control-path 
    signal convTransposeC_CP_6995_elements: BooleanArray(190 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_6995_elements(0) <= convTransposeC_CP_6995_start;
    convTransposeC_CP_6995_symbol <= convTransposeC_CP_6995_elements(141);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	45 
    -- CP-element group 0:  members (74) 
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2666/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/branch_block_stmt_2666__entry__
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970__entry__
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_Update/cr
      -- 
    cr_7734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2964_inst_req_1); -- 
    cr_7650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2926_inst_req_1); -- 
    cr_7706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2951_inst_req_1); -- 
    cr_7678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2939_inst_req_1); -- 
    rr_7043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => RPIPE_Block2_start_2668_inst_req_0); -- 
    cr_7062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2672_inst_req_1); -- 
    cr_7090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2685_inst_req_1); -- 
    cr_7118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2697_inst_req_1); -- 
    cr_7146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2710_inst_req_1); -- 
    cr_7174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2722_inst_req_1); -- 
    cr_7202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2735_inst_req_1); -- 
    cr_7258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2753_inst_req_1); -- 
    cr_7286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2766_inst_req_1); -- 
    cr_7314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2778_inst_req_1); -- 
    cr_7342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2791_inst_req_1); -- 
    cr_7398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2809_inst_req_1); -- 
    cr_7426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2822_inst_req_1); -- 
    cr_7454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2834_inst_req_1); -- 
    cr_7482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2847_inst_req_1); -- 
    cr_7510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2859_inst_req_1); -- 
    cr_7538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2872_inst_req_1); -- 
    cr_7566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2890_inst_req_1); -- 
    cr_7594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(0), ack => type_cast_2908_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	190 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	152 
    -- CP-element group 1: 	153 
    -- CP-element group 1: 	158 
    -- CP-element group 1: 	159 
    -- CP-element group 1: 	155 
    -- CP-element group 1: 	156 
    -- CP-element group 1: 	149 
    -- CP-element group 1: 	150 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2666/merge_stmt_3234__exit__
      -- CP-element group 1: 	 branch_block_stmt_2666/assign_stmt_3260__entry__
      -- CP-element group 1: 	 branch_block_stmt_2666/assign_stmt_3260__exit__
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2666/assign_stmt_3260/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/assign_stmt_3260/$exit
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/Update/cr
      -- 
    rr_8192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(1), ack => type_cast_3029_inst_req_0); -- 
    cr_8197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(1), ack => type_cast_3029_inst_req_1); -- 
    rr_8215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(1), ack => type_cast_3036_inst_req_0); -- 
    cr_8220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(1), ack => type_cast_3036_inst_req_1); -- 
    rr_8238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(1), ack => type_cast_3043_inst_req_0); -- 
    cr_8243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(1), ack => type_cast_3043_inst_req_1); -- 
    rr_8261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(1), ack => type_cast_3049_inst_req_0); -- 
    cr_8266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(1), ack => type_cast_3049_inst_req_1); -- 
    convTransposeC_CP_6995_elements(1) <= convTransposeC_CP_6995_elements(190);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_Update/cr
      -- 
    ra_7044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2668_inst_ack_0, ack => convTransposeC_CP_6995_elements(2)); -- 
    cr_7048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(2), ack => RPIPE_Block2_start_2668_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2668_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_Sample/rr
      -- 
    ca_7049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2668_inst_ack_1, ack => convTransposeC_CP_6995_elements(3)); -- 
    rr_7057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(3), ack => type_cast_2672_inst_req_0); -- 
    rr_7071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(3), ack => RPIPE_Block2_start_2681_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_Sample/ra
      -- 
    ra_7058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2672_inst_ack_0, ack => convTransposeC_CP_6995_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	102 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2672_Update/ca
      -- 
    ca_7063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2672_inst_ack_1, ack => convTransposeC_CP_6995_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_Update/cr
      -- 
    ra_7072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2681_inst_ack_0, ack => convTransposeC_CP_6995_elements(6)); -- 
    cr_7076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(6), ack => RPIPE_Block2_start_2681_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2681_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_Sample/rr
      -- 
    ca_7077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2681_inst_ack_1, ack => convTransposeC_CP_6995_elements(7)); -- 
    rr_7085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(7), ack => type_cast_2685_inst_req_0); -- 
    rr_7099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(7), ack => RPIPE_Block2_start_2693_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_Sample/ra
      -- 
    ra_7086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2685_inst_ack_0, ack => convTransposeC_CP_6995_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	102 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2685_Update/ca
      -- 
    ca_7091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2685_inst_ack_1, ack => convTransposeC_CP_6995_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_Update/cr
      -- 
    ra_7100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2693_inst_ack_0, ack => convTransposeC_CP_6995_elements(10)); -- 
    cr_7104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(10), ack => RPIPE_Block2_start_2693_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2693_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_Sample/rr
      -- 
    ca_7105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2693_inst_ack_1, ack => convTransposeC_CP_6995_elements(11)); -- 
    rr_7113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(11), ack => type_cast_2697_inst_req_0); -- 
    rr_7127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(11), ack => RPIPE_Block2_start_2706_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_Sample/ra
      -- 
    ra_7114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2697_inst_ack_0, ack => convTransposeC_CP_6995_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	102 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2697_Update/ca
      -- 
    ca_7119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2697_inst_ack_1, ack => convTransposeC_CP_6995_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_Update/cr
      -- 
    ra_7128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2706_inst_ack_0, ack => convTransposeC_CP_6995_elements(14)); -- 
    cr_7132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(14), ack => RPIPE_Block2_start_2706_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2706_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_Sample/rr
      -- 
    ca_7133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2706_inst_ack_1, ack => convTransposeC_CP_6995_elements(15)); -- 
    rr_7141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(15), ack => type_cast_2710_inst_req_0); -- 
    rr_7155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(15), ack => RPIPE_Block2_start_2718_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_Sample/ra
      -- 
    ra_7142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_0, ack => convTransposeC_CP_6995_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	102 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2710_Update/ca
      -- 
    ca_7147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2710_inst_ack_1, ack => convTransposeC_CP_6995_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_Update/cr
      -- 
    ra_7156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2718_inst_ack_0, ack => convTransposeC_CP_6995_elements(18)); -- 
    cr_7160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(18), ack => RPIPE_Block2_start_2718_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2718_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_Sample/rr
      -- 
    ca_7161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2718_inst_ack_1, ack => convTransposeC_CP_6995_elements(19)); -- 
    rr_7169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(19), ack => type_cast_2722_inst_req_0); -- 
    rr_7183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(19), ack => RPIPE_Block2_start_2731_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_Sample/ra
      -- 
    ra_7170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_0, ack => convTransposeC_CP_6995_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	102 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2722_Update/ca
      -- 
    ca_7175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_1, ack => convTransposeC_CP_6995_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_update_start_
      -- CP-element group 22: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_Update/cr
      -- 
    ra_7184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2731_inst_ack_0, ack => convTransposeC_CP_6995_elements(22)); -- 
    cr_7188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(22), ack => RPIPE_Block2_start_2731_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2731_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_Sample/rr
      -- 
    ca_7189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2731_inst_ack_1, ack => convTransposeC_CP_6995_elements(23)); -- 
    rr_7197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(23), ack => type_cast_2735_inst_req_0); -- 
    rr_7211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(23), ack => RPIPE_Block2_start_2743_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_Sample/ra
      -- 
    ra_7198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2735_inst_ack_0, ack => convTransposeC_CP_6995_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	102 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2735_Update/ca
      -- 
    ca_7203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2735_inst_ack_1, ack => convTransposeC_CP_6995_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_update_start_
      -- CP-element group 26: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_Update/cr
      -- 
    ra_7212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2743_inst_ack_0, ack => convTransposeC_CP_6995_elements(26)); -- 
    cr_7216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(26), ack => RPIPE_Block2_start_2743_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2743_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_Sample/rr
      -- 
    ca_7217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2743_inst_ack_1, ack => convTransposeC_CP_6995_elements(27)); -- 
    rr_7225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(27), ack => RPIPE_Block2_start_2746_inst_req_0); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_Update/cr
      -- 
    ra_7226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2746_inst_ack_0, ack => convTransposeC_CP_6995_elements(28)); -- 
    cr_7230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(28), ack => RPIPE_Block2_start_2746_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2746_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_Sample/rr
      -- 
    ca_7231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2746_inst_ack_1, ack => convTransposeC_CP_6995_elements(29)); -- 
    rr_7239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(29), ack => RPIPE_Block2_start_2749_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_Update/cr
      -- 
    ra_7240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2749_inst_ack_0, ack => convTransposeC_CP_6995_elements(30)); -- 
    cr_7244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(30), ack => RPIPE_Block2_start_2749_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2749_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_Sample/rr
      -- 
    ca_7245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2749_inst_ack_1, ack => convTransposeC_CP_6995_elements(31)); -- 
    rr_7253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(31), ack => type_cast_2753_inst_req_0); -- 
    rr_7267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(31), ack => RPIPE_Block2_start_2762_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_Sample/ra
      -- 
    ra_7254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2753_inst_ack_0, ack => convTransposeC_CP_6995_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	102 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2753_Update/ca
      -- 
    ca_7259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2753_inst_ack_1, ack => convTransposeC_CP_6995_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_Update/cr
      -- 
    ra_7268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2762_inst_ack_0, ack => convTransposeC_CP_6995_elements(34)); -- 
    cr_7272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(34), ack => RPIPE_Block2_start_2762_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2762_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_Sample/rr
      -- 
    ca_7273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2762_inst_ack_1, ack => convTransposeC_CP_6995_elements(35)); -- 
    rr_7281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(35), ack => type_cast_2766_inst_req_0); -- 
    rr_7295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(35), ack => RPIPE_Block2_start_2774_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_Sample/ra
      -- 
    ra_7282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_0, ack => convTransposeC_CP_6995_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	102 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2766_Update/ca
      -- 
    ca_7287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_1, ack => convTransposeC_CP_6995_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_update_start_
      -- CP-element group 38: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_Update/cr
      -- 
    ra_7296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2774_inst_ack_0, ack => convTransposeC_CP_6995_elements(38)); -- 
    cr_7300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(38), ack => RPIPE_Block2_start_2774_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2774_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_Sample/rr
      -- 
    ca_7301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2774_inst_ack_1, ack => convTransposeC_CP_6995_elements(39)); -- 
    rr_7309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(39), ack => type_cast_2778_inst_req_0); -- 
    rr_7323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(39), ack => RPIPE_Block2_start_2787_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_Sample/ra
      -- 
    ra_7310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2778_inst_ack_0, ack => convTransposeC_CP_6995_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	102 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2778_Update/ca
      -- 
    ca_7315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2778_inst_ack_1, ack => convTransposeC_CP_6995_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_update_start_
      -- CP-element group 42: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_Update/cr
      -- 
    ra_7324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2787_inst_ack_0, ack => convTransposeC_CP_6995_elements(42)); -- 
    cr_7328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(42), ack => RPIPE_Block2_start_2787_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2787_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_Sample/rr
      -- 
    ca_7329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2787_inst_ack_1, ack => convTransposeC_CP_6995_elements(43)); -- 
    rr_7337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(43), ack => type_cast_2791_inst_req_0); -- 
    rr_7351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(43), ack => RPIPE_Block2_start_2799_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_Sample/ra
      -- 
    ra_7338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2791_inst_ack_0, ack => convTransposeC_CP_6995_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	102 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2791_Update/ca
      -- 
    ca_7343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2791_inst_ack_1, ack => convTransposeC_CP_6995_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_update_start_
      -- CP-element group 46: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_Update/cr
      -- 
    ra_7352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2799_inst_ack_0, ack => convTransposeC_CP_6995_elements(46)); -- 
    cr_7356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(46), ack => RPIPE_Block2_start_2799_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2799_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_Sample/rr
      -- 
    ca_7357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2799_inst_ack_1, ack => convTransposeC_CP_6995_elements(47)); -- 
    rr_7365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(47), ack => RPIPE_Block2_start_2802_inst_req_0); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_update_start_
      -- CP-element group 48: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_Update/cr
      -- 
    ra_7366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2802_inst_ack_0, ack => convTransposeC_CP_6995_elements(48)); -- 
    cr_7370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(48), ack => RPIPE_Block2_start_2802_inst_req_1); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2802_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_Sample/rr
      -- 
    ca_7371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2802_inst_ack_1, ack => convTransposeC_CP_6995_elements(49)); -- 
    rr_7379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(49), ack => RPIPE_Block2_start_2805_inst_req_0); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_update_start_
      -- CP-element group 50: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_Update/cr
      -- 
    ra_7380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2805_inst_ack_0, ack => convTransposeC_CP_6995_elements(50)); -- 
    cr_7384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(50), ack => RPIPE_Block2_start_2805_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	54 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2805_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_Sample/rr
      -- 
    ca_7385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2805_inst_ack_1, ack => convTransposeC_CP_6995_elements(51)); -- 
    rr_7407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(51), ack => RPIPE_Block2_start_2818_inst_req_0); -- 
    rr_7393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(51), ack => type_cast_2809_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_Sample/ra
      -- 
    ra_7394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2809_inst_ack_0, ack => convTransposeC_CP_6995_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	102 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2809_Update/ca
      -- 
    ca_7399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2809_inst_ack_1, ack => convTransposeC_CP_6995_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_update_start_
      -- CP-element group 54: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_Update/cr
      -- 
    ra_7408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2818_inst_ack_0, ack => convTransposeC_CP_6995_elements(54)); -- 
    cr_7412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(54), ack => RPIPE_Block2_start_2818_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2818_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_Sample/rr
      -- 
    ca_7413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2818_inst_ack_1, ack => convTransposeC_CP_6995_elements(55)); -- 
    rr_7435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(55), ack => RPIPE_Block2_start_2830_inst_req_0); -- 
    rr_7421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(55), ack => type_cast_2822_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_Sample/ra
      -- 
    ra_7422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_0, ack => convTransposeC_CP_6995_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	102 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2822_Update/ca
      -- 
    ca_7427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2822_inst_ack_1, ack => convTransposeC_CP_6995_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_update_start_
      -- CP-element group 58: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_Update/cr
      -- 
    ra_7436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2830_inst_ack_0, ack => convTransposeC_CP_6995_elements(58)); -- 
    cr_7440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(58), ack => RPIPE_Block2_start_2830_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	62 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2830_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_Sample/rr
      -- 
    ca_7441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2830_inst_ack_1, ack => convTransposeC_CP_6995_elements(59)); -- 
    rr_7449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(59), ack => type_cast_2834_inst_req_0); -- 
    rr_7463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(59), ack => RPIPE_Block2_start_2843_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_Sample/ra
      -- 
    ra_7450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2834_inst_ack_0, ack => convTransposeC_CP_6995_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	102 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2834_Update/ca
      -- 
    ca_7455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2834_inst_ack_1, ack => convTransposeC_CP_6995_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_Update/cr
      -- 
    ra_7464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2843_inst_ack_0, ack => convTransposeC_CP_6995_elements(62)); -- 
    cr_7468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(62), ack => RPIPE_Block2_start_2843_inst_req_1); -- 
    -- CP-element group 63:  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2843_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_Sample/rr
      -- 
    ca_7469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2843_inst_ack_1, ack => convTransposeC_CP_6995_elements(63)); -- 
    rr_7477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(63), ack => type_cast_2847_inst_req_0); -- 
    rr_7491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(63), ack => RPIPE_Block2_start_2855_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_Sample/ra
      -- 
    ra_7478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2847_inst_ack_0, ack => convTransposeC_CP_6995_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	102 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2847_Update/ca
      -- 
    ca_7483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2847_inst_ack_1, ack => convTransposeC_CP_6995_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_update_start_
      -- CP-element group 66: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_Update/cr
      -- 
    ra_7492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2855_inst_ack_0, ack => convTransposeC_CP_6995_elements(66)); -- 
    cr_7496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(66), ack => RPIPE_Block2_start_2855_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	70 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2855_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_Sample/rr
      -- 
    ca_7497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2855_inst_ack_1, ack => convTransposeC_CP_6995_elements(67)); -- 
    rr_7519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(67), ack => RPIPE_Block2_start_2868_inst_req_0); -- 
    rr_7505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(67), ack => type_cast_2859_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_Sample/ra
      -- 
    ra_7506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2859_inst_ack_0, ack => convTransposeC_CP_6995_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	102 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2859_Update/ca
      -- 
    ca_7511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2859_inst_ack_1, ack => convTransposeC_CP_6995_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_Update/cr
      -- 
    ra_7520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2868_inst_ack_0, ack => convTransposeC_CP_6995_elements(70)); -- 
    cr_7524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(70), ack => RPIPE_Block2_start_2868_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	74 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2868_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_Sample/rr
      -- 
    ca_7525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2868_inst_ack_1, ack => convTransposeC_CP_6995_elements(71)); -- 
    rr_7533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(71), ack => type_cast_2872_inst_req_0); -- 
    rr_7547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(71), ack => RPIPE_Block2_start_2886_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_Sample/ra
      -- 
    ra_7534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2872_inst_ack_0, ack => convTransposeC_CP_6995_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	102 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2872_Update/ca
      -- 
    ca_7539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2872_inst_ack_1, ack => convTransposeC_CP_6995_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	71 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_update_start_
      -- CP-element group 74: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_Update/cr
      -- 
    ra_7548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2886_inst_ack_0, ack => convTransposeC_CP_6995_elements(74)); -- 
    cr_7552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(74), ack => RPIPE_Block2_start_2886_inst_req_1); -- 
    -- CP-element group 75:  fork  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (9) 
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2886_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_Sample/rr
      -- 
    ca_7553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2886_inst_ack_1, ack => convTransposeC_CP_6995_elements(75)); -- 
    rr_7561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(75), ack => type_cast_2890_inst_req_0); -- 
    rr_7575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(75), ack => RPIPE_Block2_start_2904_inst_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_Sample/ra
      -- 
    ra_7562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2890_inst_ack_0, ack => convTransposeC_CP_6995_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	102 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2890_Update/ca
      -- 
    ca_7567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2890_inst_ack_1, ack => convTransposeC_CP_6995_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_update_start_
      -- CP-element group 78: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_Update/cr
      -- 
    ra_7576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2904_inst_ack_0, ack => convTransposeC_CP_6995_elements(78)); -- 
    cr_7580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(78), ack => RPIPE_Block2_start_2904_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2904_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_Sample/rr
      -- 
    ca_7581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2904_inst_ack_1, ack => convTransposeC_CP_6995_elements(79)); -- 
    rr_7589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(79), ack => type_cast_2908_inst_req_0); -- 
    rr_7603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(79), ack => RPIPE_Block2_start_2916_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_Sample/ra
      -- 
    ra_7590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2908_inst_ack_0, ack => convTransposeC_CP_6995_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	102 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2908_Update/ca
      -- 
    ca_7595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2908_inst_ack_1, ack => convTransposeC_CP_6995_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_update_start_
      -- CP-element group 82: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_Update/cr
      -- 
    ra_7604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2916_inst_ack_0, ack => convTransposeC_CP_6995_elements(82)); -- 
    cr_7608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(82), ack => RPIPE_Block2_start_2916_inst_req_1); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2916_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_Sample/rr
      -- 
    ca_7609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2916_inst_ack_1, ack => convTransposeC_CP_6995_elements(83)); -- 
    rr_7617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(83), ack => RPIPE_Block2_start_2919_inst_req_0); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_update_start_
      -- CP-element group 84: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_Update/cr
      -- 
    ra_7618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2919_inst_ack_0, ack => convTransposeC_CP_6995_elements(84)); -- 
    cr_7622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(84), ack => RPIPE_Block2_start_2919_inst_req_1); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2919_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_Sample/rr
      -- 
    ca_7623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2919_inst_ack_1, ack => convTransposeC_CP_6995_elements(85)); -- 
    rr_7631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(85), ack => RPIPE_Block2_start_2922_inst_req_0); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_Sample/ra
      -- 
    ra_7632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2922_inst_ack_0, ack => convTransposeC_CP_6995_elements(86)); -- 
    cr_7636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(86), ack => RPIPE_Block2_start_2922_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2922_update_completed_
      -- 
    ca_7637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2922_inst_ack_1, ack => convTransposeC_CP_6995_elements(87)); -- 
    rr_7659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(87), ack => RPIPE_Block2_start_2935_inst_req_0); -- 
    rr_7645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(87), ack => type_cast_2926_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_Sample/$exit
      -- 
    ra_7646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2926_inst_ack_0, ack => convTransposeC_CP_6995_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	102 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2926_Update/ca
      -- 
    ca_7651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2926_inst_ack_1, ack => convTransposeC_CP_6995_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_update_start_
      -- CP-element group 90: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_Update/cr
      -- CP-element group 90: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_Update/$entry
      -- 
    ra_7660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2935_inst_ack_0, ack => convTransposeC_CP_6995_elements(90)); -- 
    cr_7664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(90), ack => RPIPE_Block2_start_2935_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	94 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2935_Update/$exit
      -- 
    ca_7665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2935_inst_ack_1, ack => convTransposeC_CP_6995_elements(91)); -- 
    rr_7673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(91), ack => type_cast_2939_inst_req_0); -- 
    rr_7687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(91), ack => RPIPE_Block2_start_2947_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_Sample/ra
      -- 
    ra_7674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2939_inst_ack_0, ack => convTransposeC_CP_6995_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	102 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2939_Update/$exit
      -- 
    ca_7679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2939_inst_ack_1, ack => convTransposeC_CP_6995_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_update_start_
      -- CP-element group 94: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_sample_completed_
      -- 
    ra_7688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2947_inst_ack_0, ack => convTransposeC_CP_6995_elements(94)); -- 
    cr_7692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(94), ack => RPIPE_Block2_start_2947_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2947_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_Sample/rr
      -- 
    ca_7693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2947_inst_ack_1, ack => convTransposeC_CP_6995_elements(95)); -- 
    rr_7715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(95), ack => RPIPE_Block2_start_2960_inst_req_0); -- 
    rr_7701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(95), ack => type_cast_2951_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_sample_completed_
      -- 
    ra_7702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2951_inst_ack_0, ack => convTransposeC_CP_6995_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	102 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2951_Update/ca
      -- 
    ca_7707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2951_inst_ack_1, ack => convTransposeC_CP_6995_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_Update/$entry
      -- 
    ra_7716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2960_inst_ack_0, ack => convTransposeC_CP_6995_elements(98)); -- 
    cr_7720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(98), ack => RPIPE_Block2_start_2960_inst_req_1); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/RPIPE_Block2_start_2960_update_completed_
      -- 
    ca_7721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2960_inst_ack_1, ack => convTransposeC_CP_6995_elements(99)); -- 
    rr_7729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(99), ack => type_cast_2964_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_Sample/$exit
      -- 
    ra_7730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2964_inst_ack_0, ack => convTransposeC_CP_6995_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/type_cast_2964_update_completed_
      -- 
    ca_7735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2964_inst_ack_1, ack => convTransposeC_CP_6995_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	89 
    -- CP-element group 102: 	101 
    -- CP-element group 102: 	81 
    -- CP-element group 102: 	69 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	97 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	77 
    -- CP-element group 102: 	73 
    -- CP-element group 102: 	93 
    -- CP-element group 102: 	61 
    -- CP-element group 102: 	5 
    -- CP-element group 102: 	9 
    -- CP-element group 102: 	13 
    -- CP-element group 102: 	17 
    -- CP-element group 102: 	21 
    -- CP-element group 102: 	25 
    -- CP-element group 102: 	33 
    -- CP-element group 102: 	37 
    -- CP-element group 102: 	41 
    -- CP-element group 102: 	45 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (10) 
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/$entry
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_update_start_
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970__exit__
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020__entry__
      -- CP-element group 102: 	 branch_block_stmt_2666/assign_stmt_2669_to_assign_stmt_2970/$exit
      -- 
    rr_7746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(102), ack => type_cast_3002_inst_req_0); -- 
    cr_7751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(102), ack => type_cast_3002_inst_req_1); -- 
    convTransposeC_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(89) & convTransposeC_CP_6995_elements(101) & convTransposeC_CP_6995_elements(81) & convTransposeC_CP_6995_elements(69) & convTransposeC_CP_6995_elements(57) & convTransposeC_CP_6995_elements(53) & convTransposeC_CP_6995_elements(97) & convTransposeC_CP_6995_elements(65) & convTransposeC_CP_6995_elements(77) & convTransposeC_CP_6995_elements(73) & convTransposeC_CP_6995_elements(93) & convTransposeC_CP_6995_elements(61) & convTransposeC_CP_6995_elements(5) & convTransposeC_CP_6995_elements(9) & convTransposeC_CP_6995_elements(13) & convTransposeC_CP_6995_elements(17) & convTransposeC_CP_6995_elements(21) & convTransposeC_CP_6995_elements(25) & convTransposeC_CP_6995_elements(33) & convTransposeC_CP_6995_elements(37) & convTransposeC_CP_6995_elements(41) & convTransposeC_CP_6995_elements(45);
      gj_convTransposeC_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_Sample/$exit
      -- 
    ra_7747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3002_inst_ack_0, ack => convTransposeC_CP_6995_elements(103)); -- 
    -- CP-element group 104:  fork  transition  place  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	142 
    -- CP-element group 104: 	143 
    -- CP-element group 104: 	144 
    -- CP-element group 104: 	145 
    -- CP-element group 104: 	146 
    -- CP-element group 104:  members (21) 
      -- CP-element group 104: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/$exit
      -- CP-element group 104: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020/type_cast_3002_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_2666/assign_stmt_2977_to_assign_stmt_3020__exit__
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3023/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3030/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3037/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/Update/cr
      -- 
    ca_7752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3002_inst_ack_1, ack => convTransposeC_CP_6995_elements(104)); -- 
    rr_8166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(104), ack => type_cast_3047_inst_req_0); -- 
    cr_8171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(104), ack => type_cast_3047_inst_req_1); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	167 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_sample_completed_
      -- 
    ra_7764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3084_inst_ack_0, ack => convTransposeC_CP_6995_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	167 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	119 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_Update/ca
      -- 
    ca_7769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3084_inst_ack_1, ack => convTransposeC_CP_6995_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	167 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_sample_completed_
      -- 
    ra_7778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3088_inst_ack_0, ack => convTransposeC_CP_6995_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	167 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_update_completed_
      -- 
    ca_7783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3088_inst_ack_1, ack => convTransposeC_CP_6995_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	167 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_sample_completed_
      -- 
    ra_7792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3092_inst_ack_0, ack => convTransposeC_CP_6995_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	167 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	119 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_Update/ca
      -- 
    ca_7797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3092_inst_ack_1, ack => convTransposeC_CP_6995_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	167 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_sample_completed_
      -- 
    ra_7806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3122_inst_ack_0, ack => convTransposeC_CP_6995_elements(111)); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	167 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (16) 
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_scale_1/scale_rename_req
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_scale_1/scale_rename_ack
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_resized_1
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_scaled_1
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_computed_1
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_resize_1/$entry
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_resize_1/$exit
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_resize_1/index_resize_req
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_Sample/req
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_resize_1/index_resize_ack
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_scale_1/$entry
      -- CP-element group 112: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_index_scale_1/$exit
      -- 
    ca_7811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3122_inst_ack_1, ack => convTransposeC_CP_6995_elements(112)); -- 
    req_7836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(112), ack => array_obj_ref_3128_index_offset_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	129 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_sample_complete
      -- CP-element group 113: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_Sample/ack
      -- CP-element group 113: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_Sample/$exit
      -- 
    ack_7837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3128_index_offset_ack_0, ack => convTransposeC_CP_6995_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	167 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (11) 
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_base_plus_offset/sum_rename_req
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_base_plus_offset/sum_rename_ack
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_base_plus_offset/$exit
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_base_plus_offset/$entry
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_Update/ack
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_offset_calculated
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_request/$entry
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_request/req
      -- CP-element group 114: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_root_address_calculated
      -- 
    ack_7842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3128_index_offset_ack_1, ack => convTransposeC_CP_6995_elements(114)); -- 
    req_7851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(114), ack => addr_of_3129_final_reg_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_request/$exit
      -- CP-element group 115: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_request/ack
      -- 
    ack_7852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3129_final_reg_ack_0, ack => convTransposeC_CP_6995_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	167 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (24) 
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_word_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_plus_offset/$exit
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_complete/ack
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_root_address_calculated
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_plus_offset/sum_rename_req
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_address_resized
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Sample/word_access_start/$entry
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_plus_offset/sum_rename_ack
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_addr_resize/$entry
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_word_addrgen/root_register_ack
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_complete/$exit
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_addr_resize/$exit
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_word_addrgen/$entry
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_word_addrgen/$exit
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_addr_resize/base_resize_req
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Sample/word_access_start/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_addr_resize/base_resize_ack
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_word_addrgen/root_register_req
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_base_plus_offset/$entry
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Sample/word_access_start/word_0/rr
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_update_completed_
      -- 
    ack_7857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3129_final_reg_ack_1, ack => convTransposeC_CP_6995_elements(116)); -- 
    rr_7890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(116), ack => ptr_deref_3133_load_0_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Sample/word_access_start/word_0/ra
      -- CP-element group 117: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Sample/word_access_start/word_0/$exit
      -- 
    ra_7891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3133_load_0_ack_0, ack => convTransposeC_CP_6995_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	167 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	124 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/ptr_deref_3133_Merge/$entry
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/ptr_deref_3133_Merge/$exit
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/ptr_deref_3133_Merge/merge_ack
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/ptr_deref_3133_Merge/merge_req
      -- 
    ca_7902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3133_load_0_ack_1, ack => convTransposeC_CP_6995_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	106 
    -- CP-element group 119: 	110 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (13) 
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_scaled_1
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_computed_1
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_resize_1/$entry
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_resize_1/$exit
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_resize_1/index_resize_req
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_resize_1/index_resize_ack
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_Sample/req
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_scale_1/$exit
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_resized_1
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_scale_1/scale_rename_req
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_scale_1/scale_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_index_scale_1/$entry
      -- 
    req_7932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(119), ack => array_obj_ref_3151_index_offset_req_0); -- 
    convTransposeC_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(108) & convTransposeC_CP_6995_elements(106) & convTransposeC_CP_6995_elements(110);
      gj_convTransposeC_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	129 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_Sample/ack
      -- CP-element group 120: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_sample_complete
      -- 
    ack_7933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3151_index_offset_ack_0, ack => convTransposeC_CP_6995_elements(120)); -- 
    -- CP-element group 121:  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (11) 
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_request/$entry
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_base_plus_offset/sum_rename_req
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_request/req
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_base_plus_offset/$entry
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_base_plus_offset/sum_rename_ack
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_Update/ack
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_base_plus_offset/$exit
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_root_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_offset_calculated
      -- 
    ack_7938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3151_index_offset_ack_1, ack => convTransposeC_CP_6995_elements(121)); -- 
    req_7947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(121), ack => addr_of_3152_final_reg_req_0); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_sample_completed_
      -- CP-element group 122: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_request/ack
      -- CP-element group 122: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_request/$exit
      -- 
    ack_7948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3152_final_reg_ack_0, ack => convTransposeC_CP_6995_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	167 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (19) 
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_complete/$exit
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_update_completed_
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_complete/ack
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_word_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_root_address_calculated
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_address_resized
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_addr_resize/$entry
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_addr_resize/$exit
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_addr_resize/base_resize_req
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_addr_resize/base_resize_ack
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_plus_offset/$entry
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_plus_offset/$exit
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_plus_offset/sum_rename_req
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_base_plus_offset/sum_rename_ack
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_word_addrgen/$entry
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_word_addrgen/$exit
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_word_addrgen/root_register_req
      -- CP-element group 123: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_word_addrgen/root_register_ack
      -- 
    ack_7953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3152_final_reg_ack_1, ack => convTransposeC_CP_6995_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: 	118 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/ptr_deref_3155_Split/$entry
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/ptr_deref_3155_Split/$exit
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/ptr_deref_3155_Split/split_req
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/ptr_deref_3155_Split/split_ack
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/word_access_start/$entry
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/word_access_start/word_0/$entry
      -- CP-element group 124: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/word_access_start/word_0/rr
      -- 
    rr_7991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(124), ack => ptr_deref_3155_store_0_req_0); -- 
    convTransposeC_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(123) & convTransposeC_CP_6995_elements(118);
      gj_convTransposeC_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/word_access_start/$exit
      -- CP-element group 125: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/word_access_start/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Sample/word_access_start/word_0/ra
      -- 
    ra_7992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3155_store_0_ack_0, ack => convTransposeC_CP_6995_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	167 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	129 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Update/word_access_complete/$exit
      -- CP-element group 126: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Update/word_access_complete/word_0/$exit
      -- CP-element group 126: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Update/word_access_complete/word_0/ca
      -- 
    ca_8003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3155_store_0_ack_1, ack => convTransposeC_CP_6995_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	167 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_Sample/ra
      -- 
    ra_8012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3160_inst_ack_0, ack => convTransposeC_CP_6995_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	167 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_Update/ca
      -- 
    ca_8017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3160_inst_ack_1, ack => convTransposeC_CP_6995_elements(128)); -- 
    -- CP-element group 129:  branch  join  transition  place  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	126 
    -- CP-element group 129: 	120 
    -- CP-element group 129: 	128 
    -- CP-element group 129: 	113 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (10) 
      -- CP-element group 129: 	 branch_block_stmt_2666/R_cmp_3174_place
      -- CP-element group 129: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/$exit
      -- CP-element group 129: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172__exit__
      -- CP-element group 129: 	 branch_block_stmt_2666/if_stmt_3173__entry__
      -- CP-element group 129: 	 branch_block_stmt_2666/if_stmt_3173_dead_link/$entry
      -- CP-element group 129: 	 branch_block_stmt_2666/if_stmt_3173_eval_test/$entry
      -- CP-element group 129: 	 branch_block_stmt_2666/if_stmt_3173_eval_test/$exit
      -- CP-element group 129: 	 branch_block_stmt_2666/if_stmt_3173_eval_test/branch_req
      -- CP-element group 129: 	 branch_block_stmt_2666/if_stmt_3173_if_link/$entry
      -- CP-element group 129: 	 branch_block_stmt_2666/if_stmt_3173_else_link/$entry
      -- 
    branch_req_8025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(129), ack => if_stmt_3173_branch_req_0); -- 
    convTransposeC_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(126) & convTransposeC_CP_6995_elements(120) & convTransposeC_CP_6995_elements(128) & convTransposeC_CP_6995_elements(113);
      gj_convTransposeC_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	176 
    -- CP-element group 130: 	177 
    -- CP-element group 130: 	179 
    -- CP-element group 130: 	182 
    -- CP-element group 130: 	183 
    -- CP-element group 130: 	180 
    -- CP-element group 130:  members (40) 
      -- CP-element group 130: 	 branch_block_stmt_2666/whilex_xbody_ifx_xthen
      -- CP-element group 130: 	 branch_block_stmt_2666/merge_stmt_3179__exit__
      -- CP-element group 130: 	 branch_block_stmt_2666/assign_stmt_3185__entry__
      -- CP-element group 130: 	 branch_block_stmt_2666/assign_stmt_3185__exit__
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259
      -- CP-element group 130: 	 branch_block_stmt_2666/if_stmt_3173_if_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_2666/if_stmt_3173_if_link/if_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_2666/assign_stmt_3185/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/assign_stmt_3185/$exit
      -- CP-element group 130: 	 branch_block_stmt_2666/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_2666/merge_stmt_3179_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_2666/merge_stmt_3179_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/merge_stmt_3179_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_2666/merge_stmt_3179_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/Update/cr
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/Update/cr
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/Update/cr
      -- 
    if_choice_transition_8030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3173_branch_ack_1, ack => convTransposeC_CP_6995_elements(130)); -- 
    rr_8376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(130), ack => type_cast_3238_inst_req_0); -- 
    cr_8381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(130), ack => type_cast_3238_inst_req_1); -- 
    rr_8399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(130), ack => type_cast_3245_inst_req_0); -- 
    cr_8404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(130), ack => type_cast_3245_inst_req_1); -- 
    rr_8422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(130), ack => type_cast_3251_inst_req_0); -- 
    cr_8427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(130), ack => type_cast_3251_inst_req_1); -- 
    -- CP-element group 131:  fork  transition  place  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	137 
    -- CP-element group 131: 	135 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (24) 
      -- CP-element group 131: 	 branch_block_stmt_2666/whilex_xbody_ifx_xelse
      -- CP-element group 131: 	 branch_block_stmt_2666/merge_stmt_3187__exit__
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227__entry__
      -- CP-element group 131: 	 branch_block_stmt_2666/if_stmt_3173_else_link/$exit
      -- CP-element group 131: 	 branch_block_stmt_2666/if_stmt_3173_else_link/else_choice_transition
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/$entry
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_update_start_
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_update_start_
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_update_start_
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_2666/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 131: 	 branch_block_stmt_2666/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 131: 	 branch_block_stmt_2666/merge_stmt_3187_PhiReqMerge
      -- CP-element group 131: 	 branch_block_stmt_2666/merge_stmt_3187_PhiAck/$entry
      -- CP-element group 131: 	 branch_block_stmt_2666/merge_stmt_3187_PhiAck/$exit
      -- CP-element group 131: 	 branch_block_stmt_2666/merge_stmt_3187_PhiAck/dummy
      -- 
    else_choice_transition_8034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3173_branch_ack_0, ack => convTransposeC_CP_6995_elements(131)); -- 
    rr_8050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(131), ack => type_cast_3196_inst_req_0); -- 
    cr_8055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(131), ack => type_cast_3196_inst_req_1); -- 
    cr_8069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(131), ack => type_cast_3205_inst_req_1); -- 
    cr_8083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(131), ack => type_cast_3221_inst_req_1); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_Sample/ra
      -- 
    ra_8051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3196_inst_ack_0, ack => convTransposeC_CP_6995_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3196_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_Sample/rr
      -- 
    ca_8056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3196_inst_ack_1, ack => convTransposeC_CP_6995_elements(133)); -- 
    rr_8064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(133), ack => type_cast_3205_inst_req_0); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_Sample/ra
      -- 
    ra_8065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3205_inst_ack_0, ack => convTransposeC_CP_6995_elements(134)); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	131 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (6) 
      -- CP-element group 135: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3205_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_Sample/rr
      -- 
    ca_8070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3205_inst_ack_1, ack => convTransposeC_CP_6995_elements(135)); -- 
    rr_8078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(135), ack => type_cast_3221_inst_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_Sample/ra
      -- 
    ra_8079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3221_inst_ack_0, ack => convTransposeC_CP_6995_elements(136)); -- 
    -- CP-element group 137:  branch  transition  place  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	131 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (13) 
      -- CP-element group 137: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227__exit__
      -- CP-element group 137: 	 branch_block_stmt_2666/if_stmt_3228__entry__
      -- CP-element group 137: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/$exit
      -- CP-element group 137: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_2666/assign_stmt_3193_to_assign_stmt_3227/type_cast_3221_Update/ca
      -- CP-element group 137: 	 branch_block_stmt_2666/if_stmt_3228_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_2666/if_stmt_3228_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_2666/if_stmt_3228_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_2666/if_stmt_3228_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_2666/R_cmp248_3229_place
      -- CP-element group 137: 	 branch_block_stmt_2666/if_stmt_3228_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_2666/if_stmt_3228_else_link/$entry
      -- 
    ca_8084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3221_inst_ack_1, ack => convTransposeC_CP_6995_elements(137)); -- 
    branch_req_8092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(137), ack => if_stmt_3228_branch_req_0); -- 
    -- CP-element group 138:  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (15) 
      -- CP-element group 138: 	 branch_block_stmt_2666/merge_stmt_3262__exit__
      -- CP-element group 138: 	 branch_block_stmt_2666/assign_stmt_3267__entry__
      -- CP-element group 138: 	 branch_block_stmt_2666/if_stmt_3228_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_2666/if_stmt_3228_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_2666/ifx_xelse_whilex_xend
      -- CP-element group 138: 	 branch_block_stmt_2666/assign_stmt_3267/$entry
      -- CP-element group 138: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_Sample/req
      -- CP-element group 138: 	 branch_block_stmt_2666/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_2666/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 138: 	 branch_block_stmt_2666/merge_stmt_3262_PhiReqMerge
      -- CP-element group 138: 	 branch_block_stmt_2666/merge_stmt_3262_PhiAck/$entry
      -- CP-element group 138: 	 branch_block_stmt_2666/merge_stmt_3262_PhiAck/$exit
      -- CP-element group 138: 	 branch_block_stmt_2666/merge_stmt_3262_PhiAck/dummy
      -- 
    if_choice_transition_8097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3228_branch_ack_1, ack => convTransposeC_CP_6995_elements(138)); -- 
    req_8117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(138), ack => WPIPE_Block2_done_3264_inst_req_0); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	168 
    -- CP-element group 139: 	169 
    -- CP-element group 139: 	170 
    -- CP-element group 139: 	172 
    -- CP-element group 139: 	173 
    -- CP-element group 139:  members (22) 
      -- CP-element group 139: 	 branch_block_stmt_2666/if_stmt_3228_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_2666/if_stmt_3228_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3235/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/Update/cr
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3228_branch_ack_0, ack => convTransposeC_CP_6995_elements(139)); -- 
    rr_8327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(139), ack => type_cast_3247_inst_req_0); -- 
    cr_8332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(139), ack => type_cast_3247_inst_req_1); -- 
    rr_8350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(139), ack => type_cast_3253_inst_req_0); -- 
    cr_8355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(139), ack => type_cast_3253_inst_req_1); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (6) 
      -- CP-element group 140: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_update_start_
      -- CP-element group 140: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_Sample/ack
      -- CP-element group 140: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_Update/req
      -- 
    ack_8118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_3264_inst_ack_0, ack => convTransposeC_CP_6995_elements(140)); -- 
    req_8122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(140), ack => WPIPE_Block2_done_3264_inst_req_1); -- 
    -- CP-element group 141:  transition  place  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (16) 
      -- CP-element group 141: 	 $exit
      -- CP-element group 141: 	 branch_block_stmt_2666/$exit
      -- CP-element group 141: 	 branch_block_stmt_2666/branch_block_stmt_2666__exit__
      -- CP-element group 141: 	 branch_block_stmt_2666/assign_stmt_3267__exit__
      -- CP-element group 141: 	 branch_block_stmt_2666/return__
      -- CP-element group 141: 	 branch_block_stmt_2666/merge_stmt_3269__exit__
      -- CP-element group 141: 	 branch_block_stmt_2666/assign_stmt_3267/$exit
      -- CP-element group 141: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_2666/assign_stmt_3267/WPIPE_Block2_done_3264_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_2666/return___PhiReq/$entry
      -- CP-element group 141: 	 branch_block_stmt_2666/return___PhiReq/$exit
      -- CP-element group 141: 	 branch_block_stmt_2666/merge_stmt_3269_PhiReqMerge
      -- CP-element group 141: 	 branch_block_stmt_2666/merge_stmt_3269_PhiAck/$entry
      -- CP-element group 141: 	 branch_block_stmt_2666/merge_stmt_3269_PhiAck/$exit
      -- CP-element group 141: 	 branch_block_stmt_2666/merge_stmt_3269_PhiAck/dummy
      -- 
    ack_8123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_3264_inst_ack_1, ack => convTransposeC_CP_6995_elements(141)); -- 
    -- CP-element group 142:  transition  output  delay-element  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	104 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	148 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3023/$exit
      -- CP-element group 142: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/$exit
      -- CP-element group 142: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3027_konst_delay_trans
      -- CP-element group 142: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_req
      -- 
    phi_stmt_3023_req_8134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3023_req_8134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(142), ack => phi_stmt_3023_req_0); -- 
    -- Element group convTransposeC_CP_6995_elements(142) is a control-delay.
    cp_element_142_delay: control_delay_element  generic map(name => " 142_delay", delay_value => 1)  port map(req => convTransposeC_CP_6995_elements(104), ack => convTransposeC_CP_6995_elements(142), clk => clk, reset =>reset);
    -- CP-element group 143:  transition  output  delay-element  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	104 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	148 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3030/$exit
      -- CP-element group 143: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/$exit
      -- CP-element group 143: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3034_konst_delay_trans
      -- CP-element group 143: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_req
      -- 
    phi_stmt_3030_req_8142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3030_req_8142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(143), ack => phi_stmt_3030_req_0); -- 
    -- Element group convTransposeC_CP_6995_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => convTransposeC_CP_6995_elements(104), ack => convTransposeC_CP_6995_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  transition  output  delay-element  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	104 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	148 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3037/$exit
      -- CP-element group 144: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/$exit
      -- CP-element group 144: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3041_konst_delay_trans
      -- CP-element group 144: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_req
      -- 
    phi_stmt_3037_req_8150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3037_req_8150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(144), ack => phi_stmt_3037_req_0); -- 
    -- Element group convTransposeC_CP_6995_elements(144) is a control-delay.
    cp_element_144_delay: control_delay_element  generic map(name => " 144_delay", delay_value => 1)  port map(req => convTransposeC_CP_6995_elements(104), ack => convTransposeC_CP_6995_elements(144), clk => clk, reset =>reset);
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	104 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/Sample/ra
      -- 
    ra_8167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3047_inst_ack_0, ack => convTransposeC_CP_6995_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	104 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/Update/ca
      -- 
    ca_8172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3047_inst_ack_1, ack => convTransposeC_CP_6995_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/$exit
      -- CP-element group 147: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/$exit
      -- CP-element group 147: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/$exit
      -- CP-element group 147: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3047/SplitProtocol/$exit
      -- CP-element group 147: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_req
      -- 
    phi_stmt_3044_req_8173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3044_req_8173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(147), ack => phi_stmt_3044_req_0); -- 
    convTransposeC_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(145) & convTransposeC_CP_6995_elements(146);
      gj_convTransposeC_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	142 
    -- CP-element group 148: 	143 
    -- CP-element group 148: 	144 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	162 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_2666/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(142) & convTransposeC_CP_6995_elements(143) & convTransposeC_CP_6995_elements(144) & convTransposeC_CP_6995_elements(147);
      gj_convTransposeC_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	1 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/Sample/ra
      -- 
    ra_8193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3029_inst_ack_0, ack => convTransposeC_CP_6995_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	1 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (2) 
      -- CP-element group 150: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/Update/ca
      -- 
    ca_8198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3029_inst_ack_1, ack => convTransposeC_CP_6995_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	161 
    -- CP-element group 151:  members (5) 
      -- CP-element group 151: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/$exit
      -- CP-element group 151: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/$exit
      -- CP-element group 151: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/$exit
      -- CP-element group 151: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_sources/type_cast_3029/SplitProtocol/$exit
      -- CP-element group 151: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3023/phi_stmt_3023_req
      -- 
    phi_stmt_3023_req_8199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3023_req_8199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(151), ack => phi_stmt_3023_req_1); -- 
    convTransposeC_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(149) & convTransposeC_CP_6995_elements(150);
      gj_convTransposeC_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	1 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/Sample/ra
      -- 
    ra_8216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3036_inst_ack_0, ack => convTransposeC_CP_6995_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	1 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/Update/ca
      -- 
    ca_8221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3036_inst_ack_1, ack => convTransposeC_CP_6995_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	161 
    -- CP-element group 154:  members (5) 
      -- CP-element group 154: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/$exit
      -- CP-element group 154: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/$exit
      -- CP-element group 154: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/$exit
      -- CP-element group 154: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_sources/type_cast_3036/SplitProtocol/$exit
      -- CP-element group 154: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3030/phi_stmt_3030_req
      -- 
    phi_stmt_3030_req_8222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3030_req_8222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(154), ack => phi_stmt_3030_req_1); -- 
    convTransposeC_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(152) & convTransposeC_CP_6995_elements(153);
      gj_convTransposeC_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	1 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (2) 
      -- CP-element group 155: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/Sample/ra
      -- 
    ra_8239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3043_inst_ack_0, ack => convTransposeC_CP_6995_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	1 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/Update/ca
      -- 
    ca_8244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3043_inst_ack_1, ack => convTransposeC_CP_6995_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	161 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/$exit
      -- CP-element group 157: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/$exit
      -- CP-element group 157: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/$exit
      -- CP-element group 157: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_sources/type_cast_3043/SplitProtocol/$exit
      -- CP-element group 157: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3037/phi_stmt_3037_req
      -- 
    phi_stmt_3037_req_8245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3037_req_8245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(157), ack => phi_stmt_3037_req_1); -- 
    convTransposeC_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(155) & convTransposeC_CP_6995_elements(156);
      gj_convTransposeC_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	1 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (2) 
      -- CP-element group 158: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/Sample/ra
      -- 
    ra_8262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3049_inst_ack_0, ack => convTransposeC_CP_6995_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	1 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/Update/ca
      -- 
    ca_8267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3049_inst_ack_1, ack => convTransposeC_CP_6995_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (5) 
      -- CP-element group 160: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/$exit
      -- CP-element group 160: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/$exit
      -- CP-element group 160: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/$exit
      -- CP-element group 160: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_sources/type_cast_3049/SplitProtocol/$exit
      -- CP-element group 160: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/phi_stmt_3044/phi_stmt_3044_req
      -- 
    phi_stmt_3044_req_8268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3044_req_8268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(160), ack => phi_stmt_3044_req_1); -- 
    convTransposeC_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(158) & convTransposeC_CP_6995_elements(159);
      gj_convTransposeC_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	154 
    -- CP-element group 161: 	157 
    -- CP-element group 161: 	151 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_2666/ifx_xend259_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(154) & convTransposeC_CP_6995_elements(157) & convTransposeC_CP_6995_elements(151) & convTransposeC_CP_6995_elements(160);
      gj_convTransposeC_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  merge  fork  transition  place  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	148 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	165 
    -- CP-element group 162: 	166 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (2) 
      -- CP-element group 162: 	 branch_block_stmt_2666/merge_stmt_3022_PhiReqMerge
      -- CP-element group 162: 	 branch_block_stmt_2666/merge_stmt_3022_PhiAck/$entry
      -- 
    convTransposeC_CP_6995_elements(162) <= OrReduce(convTransposeC_CP_6995_elements(148) & convTransposeC_CP_6995_elements(161));
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	167 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_2666/merge_stmt_3022_PhiAck/phi_stmt_3023_ack
      -- 
    phi_stmt_3023_ack_8273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3023_ack_0, ack => convTransposeC_CP_6995_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	167 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_2666/merge_stmt_3022_PhiAck/phi_stmt_3030_ack
      -- 
    phi_stmt_3030_ack_8274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3030_ack_0, ack => convTransposeC_CP_6995_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	162 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (1) 
      -- CP-element group 165: 	 branch_block_stmt_2666/merge_stmt_3022_PhiAck/phi_stmt_3037_ack
      -- 
    phi_stmt_3037_ack_8275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3037_ack_0, ack => convTransposeC_CP_6995_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	162 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_2666/merge_stmt_3022_PhiAck/phi_stmt_3044_ack
      -- 
    phi_stmt_3044_ack_8276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3044_ack_0, ack => convTransposeC_CP_6995_elements(166)); -- 
    -- CP-element group 167:  join  fork  transition  place  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: 	166 
    -- CP-element group 167: 	163 
    -- CP-element group 167: 	164 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	111 
    -- CP-element group 167: 	127 
    -- CP-element group 167: 	108 
    -- CP-element group 167: 	107 
    -- CP-element group 167: 	105 
    -- CP-element group 167: 	106 
    -- CP-element group 167: 	126 
    -- CP-element group 167: 	112 
    -- CP-element group 167: 	128 
    -- CP-element group 167: 	123 
    -- CP-element group 167: 	118 
    -- CP-element group 167: 	116 
    -- CP-element group 167: 	121 
    -- CP-element group 167: 	109 
    -- CP-element group 167: 	110 
    -- CP-element group 167: 	114 
    -- CP-element group 167:  members (56) 
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_update_start
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3128_final_index_sum_regn_Update/req
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_complete/req
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_Update/req
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3152_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/array_obj_ref_3151_final_index_sum_regn_update_start
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3092_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3084_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/word_access_complete/word_0/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/word_access_complete/word_0/cr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3133_Update/word_access_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3122_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/addr_of_3129_complete/req
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3088_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/merge_stmt_3022__exit__
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172__entry__
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Update/word_access_complete/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Update/word_access_complete/word_0/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/ptr_deref_3155_Update/word_access_complete/word_0/cr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_update_start_
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_2666/assign_stmt_3056_to_assign_stmt_3172/type_cast_3160_Update/cr
      -- CP-element group 167: 	 branch_block_stmt_2666/merge_stmt_3022_PhiAck/$exit
      -- 
    rr_7791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3092_inst_req_0); -- 
    rr_7805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3122_inst_req_0); -- 
    rr_7763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3084_inst_req_0); -- 
    cr_7782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3088_inst_req_1); -- 
    cr_7810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3122_inst_req_1); -- 
    rr_7777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3088_inst_req_0); -- 
    req_7841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => array_obj_ref_3128_index_offset_req_1); -- 
    req_7952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => addr_of_3152_final_reg_req_1); -- 
    req_7937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => array_obj_ref_3151_index_offset_req_1); -- 
    cr_7796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3092_inst_req_1); -- 
    cr_7768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3084_inst_req_1); -- 
    cr_7901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => ptr_deref_3133_load_0_req_1); -- 
    req_7856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => addr_of_3129_final_reg_req_1); -- 
    cr_8002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => ptr_deref_3155_store_0_req_1); -- 
    rr_8011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3160_inst_req_0); -- 
    cr_8016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(167), ack => type_cast_3160_inst_req_1); -- 
    convTransposeC_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(165) & convTransposeC_CP_6995_elements(166) & convTransposeC_CP_6995_elements(163) & convTransposeC_CP_6995_elements(164);
      gj_convTransposeC_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  transition  output  delay-element  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	139 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	175 
    -- CP-element group 168:  members (4) 
      -- CP-element group 168: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3235/$exit
      -- CP-element group 168: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/$exit
      -- CP-element group 168: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3241_konst_delay_trans
      -- CP-element group 168: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_req
      -- 
    phi_stmt_3235_req_8311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3235_req_8311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(168), ack => phi_stmt_3235_req_1); -- 
    -- Element group convTransposeC_CP_6995_elements(168) is a control-delay.
    cp_element_168_delay: control_delay_element  generic map(name => " 168_delay", delay_value => 1)  port map(req => convTransposeC_CP_6995_elements(139), ack => convTransposeC_CP_6995_elements(168), clk => clk, reset =>reset);
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	139 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (2) 
      -- CP-element group 169: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/Sample/ra
      -- 
    ra_8328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3247_inst_ack_0, ack => convTransposeC_CP_6995_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	139 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (2) 
      -- CP-element group 170: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/Update/ca
      -- 
    ca_8333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3247_inst_ack_1, ack => convTransposeC_CP_6995_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	175 
    -- CP-element group 171:  members (5) 
      -- CP-element group 171: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/$exit
      -- CP-element group 171: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/$exit
      -- CP-element group 171: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/$exit
      -- CP-element group 171: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3247/SplitProtocol/$exit
      -- CP-element group 171: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_req
      -- 
    phi_stmt_3242_req_8334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3242_req_8334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(171), ack => phi_stmt_3242_req_1); -- 
    convTransposeC_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(169) & convTransposeC_CP_6995_elements(170);
      gj_convTransposeC_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	139 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/Sample/ra
      -- 
    ra_8351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3253_inst_ack_0, ack => convTransposeC_CP_6995_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	139 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (2) 
      -- CP-element group 173: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/Update/ca
      -- 
    ca_8356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3253_inst_ack_1, ack => convTransposeC_CP_6995_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/$exit
      -- CP-element group 174: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/$exit
      -- CP-element group 174: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/$exit
      -- CP-element group 174: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3253/SplitProtocol/$exit
      -- CP-element group 174: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_req
      -- 
    phi_stmt_3248_req_8357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3248_req_8357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(174), ack => phi_stmt_3248_req_1); -- 
    convTransposeC_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(172) & convTransposeC_CP_6995_elements(173);
      gj_convTransposeC_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	171 
    -- CP-element group 175: 	168 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	186 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_2666/ifx_xelse_ifx_xend259_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(171) & convTransposeC_CP_6995_elements(168) & convTransposeC_CP_6995_elements(174);
      gj_convTransposeC_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	130 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/Sample/ra
      -- 
    ra_8377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3238_inst_ack_0, ack => convTransposeC_CP_6995_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	130 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (2) 
      -- CP-element group 177: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/Update/ca
      -- 
    ca_8382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3238_inst_ack_1, ack => convTransposeC_CP_6995_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	185 
    -- CP-element group 178:  members (5) 
      -- CP-element group 178: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/$exit
      -- CP-element group 178: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/$exit
      -- CP-element group 178: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/$exit
      -- CP-element group 178: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_sources/type_cast_3238/SplitProtocol/$exit
      -- CP-element group 178: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3235/phi_stmt_3235_req
      -- 
    phi_stmt_3235_req_8383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3235_req_8383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(178), ack => phi_stmt_3235_req_0); -- 
    convTransposeC_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(176) & convTransposeC_CP_6995_elements(177);
      gj_convTransposeC_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	130 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/Sample/ra
      -- 
    ra_8400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3245_inst_ack_0, ack => convTransposeC_CP_6995_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	130 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/Update/ca
      -- 
    ca_8405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3245_inst_ack_1, ack => convTransposeC_CP_6995_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	185 
    -- CP-element group 181:  members (5) 
      -- CP-element group 181: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/$exit
      -- CP-element group 181: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/$exit
      -- CP-element group 181: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/$exit
      -- CP-element group 181: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_sources/type_cast_3245/SplitProtocol/$exit
      -- CP-element group 181: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3242/phi_stmt_3242_req
      -- 
    phi_stmt_3242_req_8406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3242_req_8406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(181), ack => phi_stmt_3242_req_0); -- 
    convTransposeC_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(179) & convTransposeC_CP_6995_elements(180);
      gj_convTransposeC_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	130 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/Sample/ra
      -- 
    ra_8423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3251_inst_ack_0, ack => convTransposeC_CP_6995_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	130 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/Update/ca
      -- 
    ca_8428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3251_inst_ack_1, ack => convTransposeC_CP_6995_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (5) 
      -- CP-element group 184: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/$exit
      -- CP-element group 184: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/$exit
      -- CP-element group 184: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/$exit
      -- CP-element group 184: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_sources/type_cast_3251/SplitProtocol/$exit
      -- CP-element group 184: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/phi_stmt_3248/phi_stmt_3248_req
      -- 
    phi_stmt_3248_req_8429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3248_req_8429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6995_elements(184), ack => phi_stmt_3248_req_0); -- 
    convTransposeC_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(182) & convTransposeC_CP_6995_elements(183);
      gj_convTransposeC_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	178 
    -- CP-element group 185: 	181 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_2666/ifx_xthen_ifx_xend259_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(178) & convTransposeC_CP_6995_elements(181) & convTransposeC_CP_6995_elements(184);
      gj_convTransposeC_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  merge  fork  transition  place  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	175 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	189 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (2) 
      -- CP-element group 186: 	 branch_block_stmt_2666/merge_stmt_3234_PhiReqMerge
      -- CP-element group 186: 	 branch_block_stmt_2666/merge_stmt_3234_PhiAck/$entry
      -- 
    convTransposeC_CP_6995_elements(186) <= OrReduce(convTransposeC_CP_6995_elements(175) & convTransposeC_CP_6995_elements(185));
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	190 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_2666/merge_stmt_3234_PhiAck/phi_stmt_3235_ack
      -- 
    phi_stmt_3235_ack_8434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3235_ack_0, ack => convTransposeC_CP_6995_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_2666/merge_stmt_3234_PhiAck/phi_stmt_3242_ack
      -- 
    phi_stmt_3242_ack_8435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3242_ack_0, ack => convTransposeC_CP_6995_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (1) 
      -- CP-element group 189: 	 branch_block_stmt_2666/merge_stmt_3234_PhiAck/phi_stmt_3248_ack
      -- 
    phi_stmt_3248_ack_8436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3248_ack_0, ack => convTransposeC_CP_6995_elements(189)); -- 
    -- CP-element group 190:  join  transition  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: 	187 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	1 
    -- CP-element group 190:  members (1) 
      -- CP-element group 190: 	 branch_block_stmt_2666/merge_stmt_3234_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_6995_elements(189) & convTransposeC_CP_6995_elements(187) & convTransposeC_CP_6995_elements(188);
      gj_convTransposeC_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6995_elements(190), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom212_3150_resized : std_logic_vector(13 downto 0);
    signal R_idxprom212_3150_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3127_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3127_scaled : std_logic_vector(13 downto 0);
    signal add103_2878 : std_logic_vector(31 downto 0);
    signal add108_2896 : std_logic_vector(31 downto 0);
    signal add113_2914 : std_logic_vector(31 downto 0);
    signal add135_2945 : std_logic_vector(63 downto 0);
    signal add147_2970 : std_logic_vector(63 downto 0);
    signal add16_2716 : std_logic_vector(31 downto 0);
    signal add171_2983 : std_logic_vector(15 downto 0);
    signal add184_2994 : std_logic_vector(15 downto 0);
    signal add203_3103 : std_logic_vector(63 downto 0);
    signal add205_3113 : std_logic_vector(63 downto 0);
    signal add217_3167 : std_logic_vector(31 downto 0);
    signal add224_3185 : std_logic_vector(15 downto 0);
    signal add247_3020 : std_logic_vector(31 downto 0);
    signal add28_2741 : std_logic_vector(31 downto 0);
    signal add52_2772 : std_logic_vector(15 downto 0);
    signal add64_2797 : std_logic_vector(15 downto 0);
    signal add86_2828 : std_logic_vector(15 downto 0);
    signal add95_2853 : std_logic_vector(15 downto 0);
    signal add_2691 : std_logic_vector(15 downto 0);
    signal add_src_0x_x0_3061 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3128_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3128_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3128_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3128_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3128_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3128_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3151_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3151_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3151_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3151_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3151_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3151_root_address : std_logic_vector(13 downto 0);
    signal arrayidx208_3130 : std_logic_vector(31 downto 0);
    signal arrayidx213_3153 : std_logic_vector(31 downto 0);
    signal call101_2869 : std_logic_vector(7 downto 0);
    signal call106_2887 : std_logic_vector(7 downto 0);
    signal call111_2905 : std_logic_vector(7 downto 0);
    signal call114_2917 : std_logic_vector(7 downto 0);
    signal call121_2920 : std_logic_vector(7 downto 0);
    signal call126_2923 : std_logic_vector(7 downto 0);
    signal call133_2936 : std_logic_vector(7 downto 0);
    signal call138_2948 : std_logic_vector(7 downto 0);
    signal call145_2961 : std_logic_vector(7 downto 0);
    signal call14_2707 : std_logic_vector(7 downto 0);
    signal call19_2719 : std_logic_vector(7 downto 0);
    signal call26_2732 : std_logic_vector(7 downto 0);
    signal call31_2744 : std_logic_vector(7 downto 0);
    signal call38_2747 : std_logic_vector(7 downto 0);
    signal call3_2682 : std_logic_vector(7 downto 0);
    signal call43_2750 : std_logic_vector(7 downto 0);
    signal call50_2763 : std_logic_vector(7 downto 0);
    signal call55_2775 : std_logic_vector(7 downto 0);
    signal call62_2788 : std_logic_vector(7 downto 0);
    signal call67_2800 : std_logic_vector(7 downto 0);
    signal call74_2803 : std_logic_vector(7 downto 0);
    signal call79_2806 : std_logic_vector(7 downto 0);
    signal call7_2694 : std_logic_vector(7 downto 0);
    signal call84_2819 : std_logic_vector(7 downto 0);
    signal call88_2831 : std_logic_vector(7 downto 0);
    signal call93_2844 : std_logic_vector(7 downto 0);
    signal call97_2856 : std_logic_vector(7 downto 0);
    signal call_2669 : std_logic_vector(7 downto 0);
    signal cmp232_3202 : std_logic_vector(0 downto 0);
    signal cmp248_3227 : std_logic_vector(0 downto 0);
    signal cmp_3172 : std_logic_vector(0 downto 0);
    signal conv102_2873 : std_logic_vector(31 downto 0);
    signal conv107_2891 : std_logic_vector(31 downto 0);
    signal conv112_2909 : std_logic_vector(31 downto 0);
    signal conv12_2698 : std_logic_vector(31 downto 0);
    signal conv131_2927 : std_logic_vector(63 downto 0);
    signal conv134_2940 : std_logic_vector(63 downto 0);
    signal conv143_2952 : std_logic_vector(63 downto 0);
    signal conv146_2965 : std_logic_vector(63 downto 0);
    signal conv15_2711 : std_logic_vector(31 downto 0);
    signal conv191_3085 : std_logic_vector(63 downto 0);
    signal conv196_3089 : std_logic_vector(63 downto 0);
    signal conv201_3093 : std_logic_vector(63 downto 0);
    signal conv216_3161 : std_logic_vector(31 downto 0);
    signal conv228_3197 : std_logic_vector(31 downto 0);
    signal conv238_3222 : std_logic_vector(31 downto 0);
    signal conv241_3003 : std_logic_vector(31 downto 0);
    signal conv24_2723 : std_logic_vector(31 downto 0);
    signal conv27_2736 : std_logic_vector(31 downto 0);
    signal conv2_2673 : std_logic_vector(15 downto 0);
    signal conv48_2754 : std_logic_vector(15 downto 0);
    signal conv4_2686 : std_logic_vector(15 downto 0);
    signal conv51_2767 : std_logic_vector(15 downto 0);
    signal conv60_2779 : std_logic_vector(15 downto 0);
    signal conv63_2792 : std_logic_vector(15 downto 0);
    signal conv82_2810 : std_logic_vector(15 downto 0);
    signal conv85_2823 : std_logic_vector(15 downto 0);
    signal conv91_2835 : std_logic_vector(15 downto 0);
    signal conv94_2848 : std_logic_vector(15 downto 0);
    signal conv98_2860 : std_logic_vector(31 downto 0);
    signal idxprom212_3146 : std_logic_vector(63 downto 0);
    signal idxprom_3123 : std_logic_vector(63 downto 0);
    signal inc236_3206 : std_logic_vector(15 downto 0);
    signal inc236x_xinput_dim0x_x2_3211 : std_logic_vector(15 downto 0);
    signal inc_3193 : std_logic_vector(15 downto 0);
    signal indvar_3023 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_3260 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_3248 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_3044 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_3242 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_3037 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_3218 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_3235 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_3030 : std_logic_vector(15 downto 0);
    signal mul180_3076 : std_logic_vector(15 downto 0);
    signal mul202_3098 : std_logic_vector(63 downto 0);
    signal mul204_3108 : std_logic_vector(63 downto 0);
    signal mul_3066 : std_logic_vector(15 downto 0);
    signal ptr_deref_3133_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3133_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3133_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3133_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3133_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3155_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3155_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3155_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3155_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3155_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3155_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl100_2866 : std_logic_vector(31 downto 0);
    signal shl105_2884 : std_logic_vector(31 downto 0);
    signal shl110_2902 : std_logic_vector(31 downto 0);
    signal shl132_2933 : std_logic_vector(63 downto 0);
    signal shl13_2704 : std_logic_vector(31 downto 0);
    signal shl144_2958 : std_logic_vector(63 downto 0);
    signal shl25_2729 : std_logic_vector(31 downto 0);
    signal shl49_2760 : std_logic_vector(15 downto 0);
    signal shl61_2785 : std_logic_vector(15 downto 0);
    signal shl83_2816 : std_logic_vector(15 downto 0);
    signal shl92_2841 : std_logic_vector(15 downto 0);
    signal shl_2679 : std_logic_vector(15 downto 0);
    signal shr207_3119 : std_logic_vector(31 downto 0);
    signal shr211_3140 : std_logic_vector(63 downto 0);
    signal shr242263_3009 : std_logic_vector(31 downto 0);
    signal shr246264_3015 : std_logic_vector(31 downto 0);
    signal shr262_2977 : std_logic_vector(15 downto 0);
    signal sub174_3071 : std_logic_vector(15 downto 0);
    signal sub187_2999 : std_logic_vector(15 downto 0);
    signal sub188_3081 : std_logic_vector(15 downto 0);
    signal sub_2988 : std_logic_vector(15 downto 0);
    signal tmp1_3056 : std_logic_vector(31 downto 0);
    signal tmp209_3134 : std_logic_vector(63 downto 0);
    signal type_cast_2677_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2702_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2727_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2758_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2783_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2814_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2839_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2864_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2882_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2900_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2931_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2956_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2975_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2981_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2992_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3007_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3013_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3027_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3029_wire : std_logic_vector(31 downto 0);
    signal type_cast_3034_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3036_wire : std_logic_vector(15 downto 0);
    signal type_cast_3041_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3043_wire : std_logic_vector(15 downto 0);
    signal type_cast_3047_wire : std_logic_vector(15 downto 0);
    signal type_cast_3049_wire : std_logic_vector(15 downto 0);
    signal type_cast_3054_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3117_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3138_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3144_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3165_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3183_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3191_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3215_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3238_wire : std_logic_vector(15 downto 0);
    signal type_cast_3241_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3245_wire : std_logic_vector(15 downto 0);
    signal type_cast_3247_wire : std_logic_vector(15 downto 0);
    signal type_cast_3251_wire : std_logic_vector(15 downto 0);
    signal type_cast_3253_wire : std_logic_vector(15 downto 0);
    signal type_cast_3258_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3266_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_3128_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3128_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3128_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3128_resized_base_address <= "00000000000000";
    array_obj_ref_3151_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3151_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3151_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3151_resized_base_address <= "00000000000000";
    ptr_deref_3133_word_offset_0 <= "00000000000000";
    ptr_deref_3155_word_offset_0 <= "00000000000000";
    type_cast_2677_wire_constant <= "0000000000001000";
    type_cast_2702_wire_constant <= "00000000000000000000000000001000";
    type_cast_2727_wire_constant <= "00000000000000000000000000001000";
    type_cast_2758_wire_constant <= "0000000000001000";
    type_cast_2783_wire_constant <= "0000000000001000";
    type_cast_2814_wire_constant <= "0000000000001000";
    type_cast_2839_wire_constant <= "0000000000001000";
    type_cast_2864_wire_constant <= "00000000000000000000000000001000";
    type_cast_2882_wire_constant <= "00000000000000000000000000001000";
    type_cast_2900_wire_constant <= "00000000000000000000000000001000";
    type_cast_2931_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2956_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2975_wire_constant <= "0000000000000001";
    type_cast_2981_wire_constant <= "1111111111111111";
    type_cast_2992_wire_constant <= "1111111111111111";
    type_cast_3007_wire_constant <= "00000000000000000000000000000010";
    type_cast_3013_wire_constant <= "00000000000000000000000000000001";
    type_cast_3027_wire_constant <= "00000000000000000000000000000000";
    type_cast_3034_wire_constant <= "0000000000000000";
    type_cast_3041_wire_constant <= "0000000000000000";
    type_cast_3054_wire_constant <= "00000000000000000000000000000100";
    type_cast_3117_wire_constant <= "00000000000000000000000000000010";
    type_cast_3138_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_3144_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_3165_wire_constant <= "00000000000000000000000000000100";
    type_cast_3183_wire_constant <= "0000000000000100";
    type_cast_3191_wire_constant <= "0000000000000001";
    type_cast_3215_wire_constant <= "0000000000000000";
    type_cast_3241_wire_constant <= "0000000000000000";
    type_cast_3258_wire_constant <= "00000000000000000000000000000001";
    type_cast_3266_wire_constant <= "00000001";
    phi_stmt_3023: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3027_wire_constant & type_cast_3029_wire;
      req <= phi_stmt_3023_req_0 & phi_stmt_3023_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3023",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3023_ack_0,
          idata => idata,
          odata => indvar_3023,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3023
    phi_stmt_3030: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3034_wire_constant & type_cast_3036_wire;
      req <= phi_stmt_3030_req_0 & phi_stmt_3030_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3030",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3030_ack_0,
          idata => idata,
          odata => input_dim2x_x1_3030,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3030
    phi_stmt_3037: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3041_wire_constant & type_cast_3043_wire;
      req <= phi_stmt_3037_req_0 & phi_stmt_3037_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3037",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3037_ack_0,
          idata => idata,
          odata => input_dim1x_x1_3037,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3037
    phi_stmt_3044: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3047_wire & type_cast_3049_wire;
      req <= phi_stmt_3044_req_0 & phi_stmt_3044_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3044",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3044_ack_0,
          idata => idata,
          odata => input_dim0x_x2_3044,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3044
    phi_stmt_3235: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3238_wire & type_cast_3241_wire_constant;
      req <= phi_stmt_3235_req_0 & phi_stmt_3235_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3235",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3235_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_3235,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3235
    phi_stmt_3242: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3245_wire & type_cast_3247_wire;
      req <= phi_stmt_3242_req_0 & phi_stmt_3242_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3242",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3242_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_3242,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3242
    phi_stmt_3248: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3251_wire & type_cast_3253_wire;
      req <= phi_stmt_3248_req_0 & phi_stmt_3248_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3248",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3248_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_3248,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3248
    -- flow-through select operator MUX_3217_inst
    input_dim1x_x2_3218 <= type_cast_3215_wire_constant when (cmp232_3202(0) /=  '0') else inc_3193;
    addr_of_3129_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3129_final_reg_req_0;
      addr_of_3129_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3129_final_reg_req_1;
      addr_of_3129_final_reg_ack_1<= rack(0);
      addr_of_3129_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3129_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3128_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx208_3130,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3152_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3152_final_reg_req_0;
      addr_of_3152_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3152_final_reg_req_1;
      addr_of_3152_final_reg_ack_1<= rack(0);
      addr_of_3152_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3152_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3151_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx213_3153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2672_inst_req_0;
      type_cast_2672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2672_inst_req_1;
      type_cast_2672_inst_ack_1<= rack(0);
      type_cast_2672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2672_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2669,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_2673,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2685_inst_req_0;
      type_cast_2685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2685_inst_req_1;
      type_cast_2685_inst_ack_1<= rack(0);
      type_cast_2685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2682,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_2686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2697_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2697_inst_req_0;
      type_cast_2697_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2697_inst_req_1;
      type_cast_2697_inst_ack_1<= rack(0);
      type_cast_2697_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2697_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_2694,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_2698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2710_inst_req_0;
      type_cast_2710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2710_inst_req_1;
      type_cast_2710_inst_ack_1<= rack(0);
      type_cast_2710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_2707,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_2711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2722_inst_req_0;
      type_cast_2722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2722_inst_req_1;
      type_cast_2722_inst_ack_1<= rack(0);
      type_cast_2722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_2719,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_2723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2735_inst_req_0;
      type_cast_2735_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2735_inst_req_1;
      type_cast_2735_inst_ack_1<= rack(0);
      type_cast_2735_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2735_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_2732,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_2736,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2753_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2753_inst_req_0;
      type_cast_2753_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2753_inst_req_1;
      type_cast_2753_inst_ack_1<= rack(0);
      type_cast_2753_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2753_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call43_2750,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_2754,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2766_inst_req_0;
      type_cast_2766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2766_inst_req_1;
      type_cast_2766_inst_ack_1<= rack(0);
      type_cast_2766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_2763,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_2767,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2778_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2778_inst_req_0;
      type_cast_2778_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2778_inst_req_1;
      type_cast_2778_inst_ack_1<= rack(0);
      type_cast_2778_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2778_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_2775,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_2779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2791_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2791_inst_req_0;
      type_cast_2791_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2791_inst_req_1;
      type_cast_2791_inst_ack_1<= rack(0);
      type_cast_2791_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2791_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call62_2788,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_2792,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2809_inst_req_0;
      type_cast_2809_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2809_inst_req_1;
      type_cast_2809_inst_ack_1<= rack(0);
      type_cast_2809_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call79_2806,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_2810,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2822_inst_req_0;
      type_cast_2822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2822_inst_req_1;
      type_cast_2822_inst_ack_1<= rack(0);
      type_cast_2822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call84_2819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2834_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2834_inst_req_0;
      type_cast_2834_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2834_inst_req_1;
      type_cast_2834_inst_ack_1<= rack(0);
      type_cast_2834_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2834_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_2831,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_2835,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2847_inst_req_0;
      type_cast_2847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2847_inst_req_1;
      type_cast_2847_inst_ack_1<= rack(0);
      type_cast_2847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2847_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_2844,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2859_inst_req_0;
      type_cast_2859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2859_inst_req_1;
      type_cast_2859_inst_ack_1<= rack(0);
      type_cast_2859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_2856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_2860,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2872_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2872_inst_req_0;
      type_cast_2872_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2872_inst_req_1;
      type_cast_2872_inst_ack_1<= rack(0);
      type_cast_2872_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2872_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_2869,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv102_2873,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2890_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2890_inst_req_0;
      type_cast_2890_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2890_inst_req_1;
      type_cast_2890_inst_ack_1<= rack(0);
      type_cast_2890_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2890_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_2887,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_2891,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2908_inst_req_0;
      type_cast_2908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2908_inst_req_1;
      type_cast_2908_inst_ack_1<= rack(0);
      type_cast_2908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2908_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_2905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2909,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2926_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2926_inst_req_0;
      type_cast_2926_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2926_inst_req_1;
      type_cast_2926_inst_ack_1<= rack(0);
      type_cast_2926_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2926_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call126_2923,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_2927,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2939_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2939_inst_req_0;
      type_cast_2939_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2939_inst_req_1;
      type_cast_2939_inst_ack_1<= rack(0);
      type_cast_2939_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2939_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_2936,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_2940,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2951_inst_req_0;
      type_cast_2951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2951_inst_req_1;
      type_cast_2951_inst_ack_1<= rack(0);
      type_cast_2951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call138_2948,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_2952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2964_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2964_inst_req_0;
      type_cast_2964_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2964_inst_req_1;
      type_cast_2964_inst_ack_1<= rack(0);
      type_cast_2964_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2964_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_2961,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv146_2965,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3002_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3002_inst_req_0;
      type_cast_3002_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3002_inst_req_1;
      type_cast_3002_inst_ack_1<= rack(0);
      type_cast_3002_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3002_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_2691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_3003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3029_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3029_inst_req_0;
      type_cast_3029_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3029_inst_req_1;
      type_cast_3029_inst_ack_1<= rack(0);
      type_cast_3029_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3029_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_3260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3029_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3036_inst_req_0;
      type_cast_3036_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3036_inst_req_1;
      type_cast_3036_inst_ack_1<= rack(0);
      type_cast_3036_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3036_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_3235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3036_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3043_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3043_inst_req_0;
      type_cast_3043_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3043_inst_req_1;
      type_cast_3043_inst_ack_1<= rack(0);
      type_cast_3043_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3043_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_3242,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3043_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3047_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3047_inst_req_0;
      type_cast_3047_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3047_inst_req_1;
      type_cast_3047_inst_ack_1<= rack(0);
      type_cast_3047_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3047_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr262_2977,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3047_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3049_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3049_inst_req_0;
      type_cast_3049_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3049_inst_req_1;
      type_cast_3049_inst_ack_1<= rack(0);
      type_cast_3049_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3049_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_3248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3049_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3084_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3084_inst_req_0;
      type_cast_3084_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3084_inst_req_1;
      type_cast_3084_inst_ack_1<= rack(0);
      type_cast_3084_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3084_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_3030,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv191_3085,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3088_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3088_inst_req_0;
      type_cast_3088_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3088_inst_req_1;
      type_cast_3088_inst_ack_1<= rack(0);
      type_cast_3088_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3088_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub188_3081,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv196_3089,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3092_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3092_inst_req_0;
      type_cast_3092_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3092_inst_req_1;
      type_cast_3092_inst_ack_1<= rack(0);
      type_cast_3092_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3092_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub174_3071,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv201_3093,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3122_inst_req_0;
      type_cast_3122_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3122_inst_req_1;
      type_cast_3122_inst_ack_1<= rack(0);
      type_cast_3122_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3122_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr207_3119,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3123,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3160_inst_req_0;
      type_cast_3160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3160_inst_req_1;
      type_cast_3160_inst_ack_1<= rack(0);
      type_cast_3160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_3030,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv216_3161,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3196_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3196_inst_req_0;
      type_cast_3196_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3196_inst_req_1;
      type_cast_3196_inst_ack_1<= rack(0);
      type_cast_3196_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3196_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_3193,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv228_3197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3205_inst_req_0;
      type_cast_3205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3205_inst_req_1;
      type_cast_3205_inst_ack_1<= rack(0);
      type_cast_3205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp232_3202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc236_3206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3221_inst_req_0;
      type_cast_3221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3221_inst_req_1;
      type_cast_3221_inst_ack_1<= rack(0);
      type_cast_3221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc236x_xinput_dim0x_x2_3211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv238_3222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3238_inst_req_0;
      type_cast_3238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3238_inst_req_1;
      type_cast_3238_inst_ack_1<= rack(0);
      type_cast_3238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add224_3185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3238_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3245_inst_req_0;
      type_cast_3245_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3245_inst_req_1;
      type_cast_3245_inst_ack_1<= rack(0);
      type_cast_3245_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3245_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_3037,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3245_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3247_inst_req_0;
      type_cast_3247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3247_inst_req_1;
      type_cast_3247_inst_ack_1<= rack(0);
      type_cast_3247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_3218,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3247_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3251_inst_req_0;
      type_cast_3251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3251_inst_req_1;
      type_cast_3251_inst_ack_1<= rack(0);
      type_cast_3251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_3044,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3251_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3253_inst_req_0;
      type_cast_3253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3253_inst_req_1;
      type_cast_3253_inst_ack_1<= rack(0);
      type_cast_3253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc236x_xinput_dim0x_x2_3211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3253_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_3128_index_1_rename
    process(R_idxprom_3127_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3127_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3127_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3128_index_1_resize
    process(idxprom_3123) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3123;
      ov := iv(13 downto 0);
      R_idxprom_3127_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3128_root_address_inst
    process(array_obj_ref_3128_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3128_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3128_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3151_index_1_rename
    process(R_idxprom212_3150_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom212_3150_resized;
      ov(13 downto 0) := iv;
      R_idxprom212_3150_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3151_index_1_resize
    process(idxprom212_3146) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom212_3146;
      ov := iv(13 downto 0);
      R_idxprom212_3150_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3151_root_address_inst
    process(array_obj_ref_3151_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3151_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3151_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3133_addr_0
    process(ptr_deref_3133_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3133_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3133_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3133_base_resize
    process(arrayidx208_3130) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx208_3130;
      ov := iv(13 downto 0);
      ptr_deref_3133_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3133_gather_scatter
    process(ptr_deref_3133_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3133_data_0;
      ov(63 downto 0) := iv;
      tmp209_3134 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3133_root_address_inst
    process(ptr_deref_3133_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3133_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3133_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3155_addr_0
    process(ptr_deref_3155_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3155_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3155_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3155_base_resize
    process(arrayidx213_3153) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx213_3153;
      ov := iv(13 downto 0);
      ptr_deref_3155_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3155_gather_scatter
    process(tmp209_3134) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp209_3134;
      ov(63 downto 0) := iv;
      ptr_deref_3155_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3155_root_address_inst
    process(ptr_deref_3155_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3155_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3155_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3173_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_3172;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3173_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3173_branch_req_0,
          ack0 => if_stmt_3173_branch_ack_0,
          ack1 => if_stmt_3173_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3228_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp248_3227;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3228_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3228_branch_req_0,
          ack0 => if_stmt_3228_branch_ack_0,
          ack1 => if_stmt_3228_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2982_inst
    process(add52_2772) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add52_2772, type_cast_2981_wire_constant, tmp_var);
      add171_2983 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2993_inst
    process(add64_2797) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add64_2797, type_cast_2992_wire_constant, tmp_var);
      add184_2994 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3070_inst
    process(sub_2988, mul_3066) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2988, mul_3066, tmp_var);
      sub174_3071 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3080_inst
    process(sub187_2999, mul180_3076) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub187_2999, mul180_3076, tmp_var);
      sub188_3081 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3184_inst
    process(input_dim2x_x1_3030) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_3030, type_cast_3183_wire_constant, tmp_var);
      add224_3185 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3192_inst
    process(input_dim1x_x1_3037) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_3037, type_cast_3191_wire_constant, tmp_var);
      inc_3193 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3210_inst
    process(inc236_3206, input_dim0x_x2_3044) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc236_3206, input_dim0x_x2_3044, tmp_var);
      inc236x_xinput_dim0x_x2_3211 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3019_inst
    process(shr242263_3009, shr246264_3015) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr242263_3009, shr246264_3015, tmp_var);
      add247_3020 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3060_inst
    process(add113_2914, tmp1_3056) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add113_2914, tmp1_3056, tmp_var);
      add_src_0x_x0_3061 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3166_inst
    process(conv216_3161) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv216_3161, type_cast_3165_wire_constant, tmp_var);
      add217_3167 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3259_inst
    process(indvar_3023) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_3023, type_cast_3258_wire_constant, tmp_var);
      indvarx_xnext_3260 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_3102_inst
    process(mul202_3098, conv196_3089) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul202_3098, conv196_3089, tmp_var);
      add203_3103 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_3112_inst
    process(mul204_3108, conv191_3085) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul204_3108, conv191_3085, tmp_var);
      add205_3113 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_3145_inst
    process(shr211_3140) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr211_3140, type_cast_3144_wire_constant, tmp_var);
      idxprom212_3146 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3201_inst
    process(conv228_3197, add16_2716) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv228_3197, add16_2716, tmp_var);
      cmp232_3202 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3226_inst
    process(conv238_3222, add247_3020) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv238_3222, add247_3020, tmp_var);
      cmp248_3227 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2976_inst
    process(add_2691) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_2691, type_cast_2975_wire_constant, tmp_var);
      shr262_2977 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3008_inst
    process(conv241_3003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv241_3003, type_cast_3007_wire_constant, tmp_var);
      shr242263_3009 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3014_inst
    process(conv241_3003) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv241_3003, type_cast_3013_wire_constant, tmp_var);
      shr246264_3015 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3118_inst
    process(add_src_0x_x0_3061) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_3061, type_cast_3117_wire_constant, tmp_var);
      shr207_3119 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_3139_inst
    process(add205_3113) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add205_3113, type_cast_3138_wire_constant, tmp_var);
      shr211_3140 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3065_inst
    process(input_dim0x_x2_3044, add86_2828) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_3044, add86_2828, tmp_var);
      mul_3066 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3075_inst
    process(input_dim1x_x1_3037, add86_2828) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_3037, add86_2828, tmp_var);
      mul180_3076 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3055_inst
    process(indvar_3023) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_3023, type_cast_3054_wire_constant, tmp_var);
      tmp1_3056 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_3097_inst
    process(conv201_3093, add135_2945) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv201_3093, add135_2945, tmp_var);
      mul202_3098 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_3107_inst
    process(add203_3103, add147_2970) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add203_3103, add147_2970, tmp_var);
      mul204_3108 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2690_inst
    process(shl_2679, conv4_2686) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2679, conv4_2686, tmp_var);
      add_2691 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2771_inst
    process(shl49_2760, conv51_2767) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl49_2760, conv51_2767, tmp_var);
      add52_2772 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2796_inst
    process(shl61_2785, conv63_2792) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl61_2785, conv63_2792, tmp_var);
      add64_2797 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2827_inst
    process(shl83_2816, conv85_2823) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl83_2816, conv85_2823, tmp_var);
      add86_2828 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_2852_inst
    process(shl92_2841, conv94_2848) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_2841, conv94_2848, tmp_var);
      add95_2853 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2715_inst
    process(shl13_2704, conv15_2711) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl13_2704, conv15_2711, tmp_var);
      add16_2716 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2740_inst
    process(shl25_2729, conv27_2736) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl25_2729, conv27_2736, tmp_var);
      add28_2741 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2877_inst
    process(shl100_2866, conv102_2873) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_2866, conv102_2873, tmp_var);
      add103_2878 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2895_inst
    process(shl105_2884, conv107_2891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_2884, conv107_2891, tmp_var);
      add108_2896 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2913_inst
    process(shl110_2902, conv112_2909) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_2902, conv112_2909, tmp_var);
      add113_2914 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2944_inst
    process(shl132_2933, conv134_2940) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_2933, conv134_2940, tmp_var);
      add135_2945 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2969_inst
    process(shl144_2958, conv146_2965) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_2958, conv146_2965, tmp_var);
      add147_2970 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2678_inst
    process(conv2_2673) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv2_2673, type_cast_2677_wire_constant, tmp_var);
      shl_2679 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2759_inst
    process(conv48_2754) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_2754, type_cast_2758_wire_constant, tmp_var);
      shl49_2760 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2784_inst
    process(conv60_2779) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv60_2779, type_cast_2783_wire_constant, tmp_var);
      shl61_2785 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2815_inst
    process(conv82_2810) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv82_2810, type_cast_2814_wire_constant, tmp_var);
      shl83_2816 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_2840_inst
    process(conv91_2835) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_2835, type_cast_2839_wire_constant, tmp_var);
      shl92_2841 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2703_inst
    process(conv12_2698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv12_2698, type_cast_2702_wire_constant, tmp_var);
      shl13_2704 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2728_inst
    process(conv24_2723) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv24_2723, type_cast_2727_wire_constant, tmp_var);
      shl25_2729 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2865_inst
    process(conv98_2860) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv98_2860, type_cast_2864_wire_constant, tmp_var);
      shl100_2866 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2883_inst
    process(add103_2878) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add103_2878, type_cast_2882_wire_constant, tmp_var);
      shl105_2884 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2901_inst
    process(add108_2896) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_2896, type_cast_2900_wire_constant, tmp_var);
      shl110_2902 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2932_inst
    process(conv131_2927) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_2927, type_cast_2931_wire_constant, tmp_var);
      shl132_2933 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2957_inst
    process(conv143_2952) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv143_2952, type_cast_2956_wire_constant, tmp_var);
      shl144_2958 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2987_inst
    process(add171_2983, add95_2853) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add171_2983, add95_2853, tmp_var);
      sub_2988 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2998_inst
    process(add184_2994, add95_2853) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add184_2994, add95_2853, tmp_var);
      sub187_2999 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_3171_inst
    process(add217_3167, add28_2741) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add217_3167, add28_2741, tmp_var);
      cmp_3172 <= tmp_var; --
    end process;
    -- shared split operator group (53) : array_obj_ref_3128_index_offset 
    ApIntAdd_group_53: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3127_scaled;
      array_obj_ref_3128_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3128_index_offset_req_0;
      array_obj_ref_3128_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3128_index_offset_req_1;
      array_obj_ref_3128_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_53_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_53_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : array_obj_ref_3151_index_offset 
    ApIntAdd_group_54: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom212_3150_scaled;
      array_obj_ref_3151_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3151_index_offset_req_0;
      array_obj_ref_3151_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3151_index_offset_req_1;
      array_obj_ref_3151_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_54_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_54_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_54",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared load operator group (0) : ptr_deref_3133_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3133_load_0_req_0;
      ptr_deref_3133_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3133_load_0_req_1;
      ptr_deref_3133_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3133_word_address_0;
      ptr_deref_3133_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3155_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3155_store_0_req_0;
      ptr_deref_3155_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3155_store_0_req_1;
      ptr_deref_3155_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3155_word_address_0;
      data_in <= ptr_deref_3155_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2916_inst RPIPE_Block2_start_2868_inst RPIPE_Block2_start_2935_inst RPIPE_Block2_start_2947_inst RPIPE_Block2_start_2919_inst RPIPE_Block2_start_2922_inst RPIPE_Block2_start_2843_inst RPIPE_Block2_start_2886_inst RPIPE_Block2_start_2960_inst RPIPE_Block2_start_2904_inst RPIPE_Block2_start_2855_inst RPIPE_Block2_start_2668_inst RPIPE_Block2_start_2681_inst RPIPE_Block2_start_2693_inst RPIPE_Block2_start_2706_inst RPIPE_Block2_start_2718_inst RPIPE_Block2_start_2731_inst RPIPE_Block2_start_2743_inst RPIPE_Block2_start_2746_inst RPIPE_Block2_start_2749_inst RPIPE_Block2_start_2762_inst RPIPE_Block2_start_2774_inst RPIPE_Block2_start_2787_inst RPIPE_Block2_start_2799_inst RPIPE_Block2_start_2802_inst RPIPE_Block2_start_2805_inst RPIPE_Block2_start_2818_inst RPIPE_Block2_start_2830_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 27 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 27 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant outBUFs : IntegerArray(27 downto 0) := (27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      reqL_unguarded(27) <= RPIPE_Block2_start_2916_inst_req_0;
      reqL_unguarded(26) <= RPIPE_Block2_start_2868_inst_req_0;
      reqL_unguarded(25) <= RPIPE_Block2_start_2935_inst_req_0;
      reqL_unguarded(24) <= RPIPE_Block2_start_2947_inst_req_0;
      reqL_unguarded(23) <= RPIPE_Block2_start_2919_inst_req_0;
      reqL_unguarded(22) <= RPIPE_Block2_start_2922_inst_req_0;
      reqL_unguarded(21) <= RPIPE_Block2_start_2843_inst_req_0;
      reqL_unguarded(20) <= RPIPE_Block2_start_2886_inst_req_0;
      reqL_unguarded(19) <= RPIPE_Block2_start_2960_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Block2_start_2904_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Block2_start_2855_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Block2_start_2668_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Block2_start_2681_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Block2_start_2693_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Block2_start_2706_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2718_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2731_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2743_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2746_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2749_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2762_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2774_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2787_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2799_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2802_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2805_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2818_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2830_inst_req_0;
      RPIPE_Block2_start_2916_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_Block2_start_2868_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_Block2_start_2935_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_Block2_start_2947_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_Block2_start_2919_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_Block2_start_2922_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_Block2_start_2843_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_Block2_start_2886_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_Block2_start_2960_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Block2_start_2904_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Block2_start_2855_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Block2_start_2668_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Block2_start_2681_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Block2_start_2693_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Block2_start_2706_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2718_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2731_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2743_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2746_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2749_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2762_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2774_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2787_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2799_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2802_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2805_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2818_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2830_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(27) <= RPIPE_Block2_start_2916_inst_req_1;
      reqR_unguarded(26) <= RPIPE_Block2_start_2868_inst_req_1;
      reqR_unguarded(25) <= RPIPE_Block2_start_2935_inst_req_1;
      reqR_unguarded(24) <= RPIPE_Block2_start_2947_inst_req_1;
      reqR_unguarded(23) <= RPIPE_Block2_start_2919_inst_req_1;
      reqR_unguarded(22) <= RPIPE_Block2_start_2922_inst_req_1;
      reqR_unguarded(21) <= RPIPE_Block2_start_2843_inst_req_1;
      reqR_unguarded(20) <= RPIPE_Block2_start_2886_inst_req_1;
      reqR_unguarded(19) <= RPIPE_Block2_start_2960_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Block2_start_2904_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Block2_start_2855_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Block2_start_2668_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Block2_start_2681_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Block2_start_2693_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Block2_start_2706_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2718_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2731_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2743_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2746_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2749_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2762_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2774_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2787_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2799_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2802_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2805_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2818_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2830_inst_req_1;
      RPIPE_Block2_start_2916_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_Block2_start_2868_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_Block2_start_2935_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_Block2_start_2947_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_Block2_start_2919_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_Block2_start_2922_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_Block2_start_2843_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_Block2_start_2886_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_Block2_start_2960_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Block2_start_2904_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Block2_start_2855_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Block2_start_2668_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Block2_start_2681_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Block2_start_2693_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Block2_start_2706_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2718_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2731_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2743_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2746_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2749_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2762_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2774_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2787_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2799_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2802_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2805_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2818_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2830_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      call114_2917 <= data_out(223 downto 216);
      call101_2869 <= data_out(215 downto 208);
      call133_2936 <= data_out(207 downto 200);
      call138_2948 <= data_out(199 downto 192);
      call121_2920 <= data_out(191 downto 184);
      call126_2923 <= data_out(183 downto 176);
      call93_2844 <= data_out(175 downto 168);
      call106_2887 <= data_out(167 downto 160);
      call145_2961 <= data_out(159 downto 152);
      call111_2905 <= data_out(151 downto 144);
      call97_2856 <= data_out(143 downto 136);
      call_2669 <= data_out(135 downto 128);
      call3_2682 <= data_out(127 downto 120);
      call7_2694 <= data_out(119 downto 112);
      call14_2707 <= data_out(111 downto 104);
      call19_2719 <= data_out(103 downto 96);
      call26_2732 <= data_out(95 downto 88);
      call31_2744 <= data_out(87 downto 80);
      call38_2747 <= data_out(79 downto 72);
      call43_2750 <= data_out(71 downto 64);
      call50_2763 <= data_out(63 downto 56);
      call55_2775 <= data_out(55 downto 48);
      call62_2788 <= data_out(47 downto 40);
      call67_2800 <= data_out(39 downto 32);
      call74_2803 <= data_out(31 downto 24);
      call79_2806 <= data_out(23 downto 16);
      call84_2819 <= data_out(15 downto 8);
      call88_2831 <= data_out(7 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 8,  num_reqs => 28,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_3264_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_3264_inst_req_0;
      WPIPE_Block2_done_3264_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_3264_inst_req_1;
      WPIPE_Block2_done_3264_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_3266_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_8453_start: Boolean;
  signal convTransposeD_CP_8453_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_3304_inst_ack_0 : boolean;
  signal type_cast_3304_inst_req_1 : boolean;
  signal type_cast_3292_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3288_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3275_inst_req_0 : boolean;
  signal type_cast_3279_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3288_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3275_inst_ack_0 : boolean;
  signal type_cast_3279_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3288_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3313_inst_ack_1 : boolean;
  signal type_cast_3292_inst_ack_0 : boolean;
  signal type_cast_3685_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3275_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3288_inst_ack_1 : boolean;
  signal type_cast_3279_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3313_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3529_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3275_inst_ack_1 : boolean;
  signal type_cast_3304_inst_req_0 : boolean;
  signal type_cast_3279_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3313_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3300_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3300_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3325_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3300_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3325_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3325_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3554_inst_req_0 : boolean;
  signal type_cast_3681_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3300_inst_ack_0 : boolean;
  signal ptr_deref_3730_load_0_req_0 : boolean;
  signal RPIPE_Block3_start_3325_inst_ack_1 : boolean;
  signal ptr_deref_3730_load_0_ack_0 : boolean;
  signal addr_of_3726_final_reg_ack_0 : boolean;
  signal type_cast_3681_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3313_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3338_inst_ack_0 : boolean;
  signal type_cast_3681_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3338_inst_req_0 : boolean;
  signal type_cast_3681_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3350_inst_ack_0 : boolean;
  signal type_cast_3329_inst_ack_1 : boolean;
  signal type_cast_3317_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3350_inst_req_0 : boolean;
  signal type_cast_3329_inst_req_1 : boolean;
  signal ptr_deref_3752_store_0_req_0 : boolean;
  signal type_cast_3317_inst_req_1 : boolean;
  signal type_cast_3342_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3353_inst_ack_1 : boolean;
  signal type_cast_3342_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3353_inst_req_1 : boolean;
  signal type_cast_3329_inst_ack_0 : boolean;
  signal type_cast_3342_inst_req_0 : boolean;
  signal type_cast_3342_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3353_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3353_inst_ack_0 : boolean;
  signal type_cast_3329_inst_req_0 : boolean;
  signal type_cast_3317_inst_ack_0 : boolean;
  signal type_cast_3317_inst_req_0 : boolean;
  signal type_cast_3292_inst_ack_1 : boolean;
  signal addr_of_3749_final_reg_ack_1 : boolean;
  signal addr_of_3749_final_reg_req_1 : boolean;
  signal RPIPE_Block3_start_3529_inst_req_1 : boolean;
  signal ptr_deref_3752_store_0_ack_0 : boolean;
  signal RPIPE_Block3_start_3338_inst_ack_1 : boolean;
  signal type_cast_3292_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3350_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3350_inst_ack_1 : boolean;
  signal type_cast_3304_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3338_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3356_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3356_inst_ack_0 : boolean;
  signal type_cast_3546_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3356_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3356_inst_ack_1 : boolean;
  signal type_cast_3533_inst_ack_1 : boolean;
  signal type_cast_3533_inst_req_1 : boolean;
  signal type_cast_3533_inst_ack_0 : boolean;
  signal type_cast_3360_inst_req_0 : boolean;
  signal type_cast_3360_inst_ack_0 : boolean;
  signal type_cast_3360_inst_req_1 : boolean;
  signal type_cast_3360_inst_ack_1 : boolean;
  signal type_cast_3533_inst_req_0 : boolean;
  signal type_cast_3571_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3369_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3369_inst_ack_0 : boolean;
  signal type_cast_3546_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3369_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3369_inst_ack_1 : boolean;
  signal addr_of_3749_final_reg_ack_0 : boolean;
  signal addr_of_3749_final_reg_req_0 : boolean;
  signal type_cast_3571_inst_req_1 : boolean;
  signal type_cast_3373_inst_req_0 : boolean;
  signal type_cast_3373_inst_ack_0 : boolean;
  signal type_cast_3373_inst_req_1 : boolean;
  signal type_cast_3373_inst_ack_1 : boolean;
  signal type_cast_3571_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3381_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3381_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3381_inst_req_1 : boolean;
  signal type_cast_3719_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3381_inst_ack_1 : boolean;
  signal type_cast_3571_inst_req_0 : boolean;
  signal addr_of_3726_final_reg_ack_1 : boolean;
  signal type_cast_3385_inst_req_0 : boolean;
  signal type_cast_3719_inst_req_1 : boolean;
  signal type_cast_3385_inst_ack_0 : boolean;
  signal type_cast_3385_inst_req_1 : boolean;
  signal type_cast_3385_inst_ack_1 : boolean;
  signal addr_of_3726_final_reg_req_1 : boolean;
  signal RPIPE_Block3_start_3394_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3394_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3394_inst_req_1 : boolean;
  signal type_cast_3719_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3394_inst_ack_1 : boolean;
  signal array_obj_ref_3748_index_offset_ack_1 : boolean;
  signal ptr_deref_3752_store_0_req_1 : boolean;
  signal ptr_deref_3752_store_0_ack_1 : boolean;
  signal type_cast_3719_inst_req_0 : boolean;
  signal type_cast_3398_inst_req_0 : boolean;
  signal type_cast_3398_inst_ack_0 : boolean;
  signal type_cast_3398_inst_req_1 : boolean;
  signal type_cast_3398_inst_ack_1 : boolean;
  signal addr_of_3726_final_reg_req_0 : boolean;
  signal type_cast_3546_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3406_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3406_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3406_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3406_inst_ack_1 : boolean;
  signal array_obj_ref_3748_index_offset_req_1 : boolean;
  signal RPIPE_Block3_start_3567_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3409_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3409_inst_ack_0 : boolean;
  signal type_cast_3546_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3409_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3409_inst_ack_1 : boolean;
  signal array_obj_ref_3748_index_offset_ack_0 : boolean;
  signal array_obj_ref_3748_index_offset_req_0 : boolean;
  signal RPIPE_Block3_start_3567_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3412_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3412_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3412_inst_req_1 : boolean;
  signal type_cast_3689_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3412_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3567_inst_ack_0 : boolean;
  signal type_cast_3416_inst_req_0 : boolean;
  signal type_cast_3689_inst_req_1 : boolean;
  signal type_cast_3416_inst_ack_0 : boolean;
  signal type_cast_3416_inst_req_1 : boolean;
  signal type_cast_3416_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3567_inst_req_0 : boolean;
  signal array_obj_ref_3725_index_offset_ack_1 : boolean;
  signal RPIPE_Block3_start_3425_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3425_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3425_inst_req_1 : boolean;
  signal type_cast_3689_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3425_inst_ack_1 : boolean;
  signal type_cast_3429_inst_req_0 : boolean;
  signal type_cast_3689_inst_req_0 : boolean;
  signal type_cast_3429_inst_ack_0 : boolean;
  signal ptr_deref_3730_load_0_ack_1 : boolean;
  signal type_cast_3429_inst_req_1 : boolean;
  signal type_cast_3429_inst_ack_1 : boolean;
  signal array_obj_ref_3725_index_offset_req_1 : boolean;
  signal type_cast_3558_inst_ack_1 : boolean;
  signal type_cast_3558_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3437_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3437_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3437_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3437_inst_ack_1 : boolean;
  signal type_cast_3558_inst_ack_0 : boolean;
  signal type_cast_3558_inst_req_0 : boolean;
  signal ptr_deref_3730_load_0_req_1 : boolean;
  signal type_cast_3441_inst_req_0 : boolean;
  signal type_cast_3441_inst_ack_0 : boolean;
  signal type_cast_3441_inst_req_1 : boolean;
  signal type_cast_3441_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3542_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3542_inst_req_1 : boolean;
  signal array_obj_ref_3725_index_offset_ack_0 : boolean;
  signal RPIPE_Block3_start_3450_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3450_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3450_inst_req_1 : boolean;
  signal type_cast_3685_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3450_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3554_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3554_inst_req_1 : boolean;
  signal type_cast_3454_inst_req_0 : boolean;
  signal type_cast_3685_inst_req_1 : boolean;
  signal type_cast_3454_inst_ack_0 : boolean;
  signal type_cast_3454_inst_req_1 : boolean;
  signal type_cast_3454_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3542_inst_ack_0 : boolean;
  signal array_obj_ref_3725_index_offset_req_0 : boolean;
  signal RPIPE_Block3_start_3542_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3554_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3462_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3462_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3462_inst_req_1 : boolean;
  signal type_cast_3685_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3462_inst_ack_1 : boolean;
  signal type_cast_3466_inst_req_0 : boolean;
  signal type_cast_3466_inst_ack_0 : boolean;
  signal type_cast_3466_inst_req_1 : boolean;
  signal type_cast_3466_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3475_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3475_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3475_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3475_inst_ack_1 : boolean;
  signal type_cast_3479_inst_req_0 : boolean;
  signal type_cast_3479_inst_ack_0 : boolean;
  signal type_cast_3479_inst_req_1 : boolean;
  signal type_cast_3479_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3493_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3493_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3493_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3493_inst_ack_1 : boolean;
  signal type_cast_3497_inst_req_0 : boolean;
  signal type_cast_3497_inst_ack_0 : boolean;
  signal type_cast_3497_inst_req_1 : boolean;
  signal type_cast_3497_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3511_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3511_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3511_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3511_inst_ack_1 : boolean;
  signal type_cast_3515_inst_req_0 : boolean;
  signal type_cast_3515_inst_ack_0 : boolean;
  signal type_cast_3515_inst_req_1 : boolean;
  signal type_cast_3515_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3523_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3523_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3523_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3523_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3526_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3526_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_3526_inst_req_1 : boolean;
  signal RPIPE_Block3_start_3526_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_3529_inst_req_0 : boolean;
  signal RPIPE_Block3_start_3529_inst_ack_0 : boolean;
  signal type_cast_3757_inst_req_0 : boolean;
  signal type_cast_3757_inst_ack_0 : boolean;
  signal type_cast_3757_inst_req_1 : boolean;
  signal type_cast_3757_inst_ack_1 : boolean;
  signal if_stmt_3770_branch_req_0 : boolean;
  signal if_stmt_3770_branch_ack_1 : boolean;
  signal if_stmt_3770_branch_ack_0 : boolean;
  signal type_cast_3793_inst_req_0 : boolean;
  signal type_cast_3793_inst_ack_0 : boolean;
  signal type_cast_3793_inst_req_1 : boolean;
  signal type_cast_3793_inst_ack_1 : boolean;
  signal type_cast_3802_inst_req_0 : boolean;
  signal type_cast_3802_inst_ack_0 : boolean;
  signal type_cast_3802_inst_req_1 : boolean;
  signal type_cast_3802_inst_ack_1 : boolean;
  signal if_stmt_3821_branch_req_0 : boolean;
  signal if_stmt_3821_branch_ack_1 : boolean;
  signal if_stmt_3821_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_3857_inst_req_0 : boolean;
  signal WPIPE_Block3_done_3857_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_3857_inst_req_1 : boolean;
  signal WPIPE_Block3_done_3857_inst_ack_1 : boolean;
  signal type_cast_3646_inst_req_0 : boolean;
  signal type_cast_3646_inst_ack_0 : boolean;
  signal type_cast_3646_inst_req_1 : boolean;
  signal type_cast_3646_inst_ack_1 : boolean;
  signal phi_stmt_3641_req_1 : boolean;
  signal phi_stmt_3634_req_0 : boolean;
  signal phi_stmt_3627_req_0 : boolean;
  signal phi_stmt_3620_req_0 : boolean;
  signal type_cast_3644_inst_req_0 : boolean;
  signal type_cast_3644_inst_ack_0 : boolean;
  signal type_cast_3644_inst_req_1 : boolean;
  signal type_cast_3644_inst_ack_1 : boolean;
  signal phi_stmt_3641_req_0 : boolean;
  signal type_cast_3640_inst_req_0 : boolean;
  signal type_cast_3640_inst_ack_0 : boolean;
  signal type_cast_3640_inst_req_1 : boolean;
  signal type_cast_3640_inst_ack_1 : boolean;
  signal phi_stmt_3634_req_1 : boolean;
  signal type_cast_3633_inst_req_0 : boolean;
  signal type_cast_3633_inst_ack_0 : boolean;
  signal type_cast_3633_inst_req_1 : boolean;
  signal type_cast_3633_inst_ack_1 : boolean;
  signal phi_stmt_3627_req_1 : boolean;
  signal type_cast_3626_inst_req_0 : boolean;
  signal type_cast_3626_inst_ack_0 : boolean;
  signal type_cast_3626_inst_req_1 : boolean;
  signal type_cast_3626_inst_ack_1 : boolean;
  signal phi_stmt_3620_req_1 : boolean;
  signal phi_stmt_3620_ack_0 : boolean;
  signal phi_stmt_3627_ack_0 : boolean;
  signal phi_stmt_3634_ack_0 : boolean;
  signal phi_stmt_3641_ack_0 : boolean;
  signal type_cast_3846_inst_req_0 : boolean;
  signal type_cast_3846_inst_ack_0 : boolean;
  signal type_cast_3846_inst_req_1 : boolean;
  signal type_cast_3846_inst_ack_1 : boolean;
  signal phi_stmt_3841_req_1 : boolean;
  signal type_cast_3840_inst_req_0 : boolean;
  signal type_cast_3840_inst_ack_0 : boolean;
  signal type_cast_3840_inst_req_1 : boolean;
  signal type_cast_3840_inst_ack_1 : boolean;
  signal phi_stmt_3835_req_1 : boolean;
  signal phi_stmt_3828_req_0 : boolean;
  signal type_cast_3844_inst_req_0 : boolean;
  signal type_cast_3844_inst_ack_0 : boolean;
  signal type_cast_3844_inst_req_1 : boolean;
  signal type_cast_3844_inst_ack_1 : boolean;
  signal phi_stmt_3841_req_0 : boolean;
  signal type_cast_3838_inst_req_0 : boolean;
  signal type_cast_3838_inst_ack_0 : boolean;
  signal type_cast_3838_inst_req_1 : boolean;
  signal type_cast_3838_inst_ack_1 : boolean;
  signal phi_stmt_3835_req_0 : boolean;
  signal type_cast_3834_inst_req_0 : boolean;
  signal type_cast_3834_inst_ack_0 : boolean;
  signal type_cast_3834_inst_req_1 : boolean;
  signal type_cast_3834_inst_ack_1 : boolean;
  signal phi_stmt_3828_req_1 : boolean;
  signal phi_stmt_3828_ack_0 : boolean;
  signal phi_stmt_3835_ack_0 : boolean;
  signal phi_stmt_3841_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_8453_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_8453_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_8453_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_8453_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_8453: Block -- control-path 
    signal convTransposeD_CP_8453_elements: BooleanArray(186 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_8453_elements(0) <= convTransposeD_CP_8453_start;
    convTransposeD_CP_8453_symbol <= convTransposeD_CP_8453_elements(137);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	57 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	61 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	53 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0:  members (74) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577__entry__
      -- CP-element group 0: 	 branch_block_stmt_3273/branch_block_stmt_3273__entry__
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_update_start_
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_Update/cr
      -- 
    cr_8576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3304_inst_req_1); -- 
    rr_8501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => RPIPE_Block3_start_3275_inst_req_0); -- 
    cr_8520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3279_inst_req_1); -- 
    cr_8632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3329_inst_req_1); -- 
    cr_8604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3317_inst_req_1); -- 
    cr_8660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3342_inst_req_1); -- 
    cr_8548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3292_inst_req_1); -- 
    cr_9108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3533_inst_req_1); -- 
    cr_8716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3360_inst_req_1); -- 
    cr_9136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3546_inst_req_1); -- 
    cr_9192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3571_inst_req_1); -- 
    cr_8744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3373_inst_req_1); -- 
    cr_8772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3385_inst_req_1); -- 
    cr_8800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3398_inst_req_1); -- 
    cr_8856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3416_inst_req_1); -- 
    cr_8884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3429_inst_req_1); -- 
    cr_9164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3558_inst_req_1); -- 
    cr_8912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3441_inst_req_1); -- 
    cr_8940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3454_inst_req_1); -- 
    cr_8968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3466_inst_req_1); -- 
    cr_8996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3479_inst_req_1); -- 
    cr_9024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3497_inst_req_1); -- 
    cr_9052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(0), ack => type_cast_3515_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	186 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	148 
    -- CP-element group 1: 	149 
    -- CP-element group 1: 	154 
    -- CP-element group 1: 	155 
    -- CP-element group 1: 	151 
    -- CP-element group 1: 	152 
    -- CP-element group 1: 	145 
    -- CP-element group 1: 	146 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_3273/merge_stmt_3827__exit__
      -- CP-element group 1: 	 branch_block_stmt_3273/assign_stmt_3853__entry__
      -- CP-element group 1: 	 branch_block_stmt_3273/assign_stmt_3853__exit__
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_3273/assign_stmt_3853/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/assign_stmt_3853/$exit
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/Update/cr
      -- 
    rr_9622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(1), ack => type_cast_3644_inst_req_0); -- 
    cr_9627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(1), ack => type_cast_3644_inst_req_1); -- 
    rr_9645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(1), ack => type_cast_3640_inst_req_0); -- 
    cr_9650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(1), ack => type_cast_3640_inst_req_1); -- 
    rr_9668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(1), ack => type_cast_3633_inst_req_0); -- 
    cr_9673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(1), ack => type_cast_3633_inst_req_1); -- 
    rr_9691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(1), ack => type_cast_3626_inst_req_0); -- 
    cr_9696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(1), ack => type_cast_3626_inst_req_1); -- 
    convTransposeD_CP_8453_elements(1) <= convTransposeD_CP_8453_elements(186);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_update_start_
      -- CP-element group 2: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_Update/cr
      -- 
    ra_8502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3275_inst_ack_0, ack => convTransposeD_CP_8453_elements(2)); -- 
    cr_8506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(2), ack => RPIPE_Block3_start_3275_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3275_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_sample_start_
      -- 
    ca_8507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3275_inst_ack_1, ack => convTransposeD_CP_8453_elements(3)); -- 
    rr_8515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(3), ack => type_cast_3279_inst_req_0); -- 
    rr_8529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(3), ack => RPIPE_Block3_start_3288_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_sample_completed_
      -- 
    ra_8516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3279_inst_ack_0, ack => convTransposeD_CP_8453_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	102 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3279_update_completed_
      -- 
    ca_8521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3279_inst_ack_1, ack => convTransposeD_CP_8453_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_update_start_
      -- CP-element group 6: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_Update/cr
      -- 
    ra_8530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3288_inst_ack_0, ack => convTransposeD_CP_8453_elements(6)); -- 
    cr_8534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(6), ack => RPIPE_Block3_start_3288_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3288_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_Sample/rr
      -- 
    ca_8535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3288_inst_ack_1, ack => convTransposeD_CP_8453_elements(7)); -- 
    rr_8543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(7), ack => type_cast_3292_inst_req_0); -- 
    rr_8557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(7), ack => RPIPE_Block3_start_3300_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_sample_completed_
      -- 
    ra_8544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3292_inst_ack_0, ack => convTransposeD_CP_8453_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	102 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3292_Update/ca
      -- 
    ca_8549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3292_inst_ack_1, ack => convTransposeD_CP_8453_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_update_start_
      -- CP-element group 10: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_Sample/ra
      -- 
    ra_8558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3300_inst_ack_0, ack => convTransposeD_CP_8453_elements(10)); -- 
    cr_8562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(10), ack => RPIPE_Block3_start_3300_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3300_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_sample_start_
      -- 
    ca_8563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3300_inst_ack_1, ack => convTransposeD_CP_8453_elements(11)); -- 
    rr_8571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(11), ack => type_cast_3304_inst_req_0); -- 
    rr_8585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(11), ack => RPIPE_Block3_start_3313_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_sample_completed_
      -- 
    ra_8572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3304_inst_ack_0, ack => convTransposeD_CP_8453_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	102 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3304_Update/ca
      -- 
    ca_8577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3304_inst_ack_1, ack => convTransposeD_CP_8453_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_update_start_
      -- CP-element group 14: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_Update/cr
      -- 
    ra_8586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3313_inst_ack_0, ack => convTransposeD_CP_8453_elements(14)); -- 
    cr_8590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(14), ack => RPIPE_Block3_start_3313_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3313_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_Sample/$entry
      -- 
    ca_8591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3313_inst_ack_1, ack => convTransposeD_CP_8453_elements(15)); -- 
    rr_8599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(15), ack => type_cast_3317_inst_req_0); -- 
    rr_8613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(15), ack => RPIPE_Block3_start_3325_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_Sample/$exit
      -- 
    ra_8600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3317_inst_ack_0, ack => convTransposeD_CP_8453_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	102 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3317_Update/$exit
      -- 
    ca_8605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3317_inst_ack_1, ack => convTransposeD_CP_8453_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_update_start_
      -- CP-element group 18: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_sample_completed_
      -- 
    ra_8614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3325_inst_ack_0, ack => convTransposeD_CP_8453_elements(18)); -- 
    cr_8618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(18), ack => RPIPE_Block3_start_3325_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3325_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_sample_start_
      -- 
    ca_8619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3325_inst_ack_1, ack => convTransposeD_CP_8453_elements(19)); -- 
    rr_8627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(19), ack => type_cast_3329_inst_req_0); -- 
    rr_8641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(19), ack => RPIPE_Block3_start_3338_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_sample_completed_
      -- 
    ra_8628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3329_inst_ack_0, ack => convTransposeD_CP_8453_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	102 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3329_update_completed_
      -- 
    ca_8633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3329_inst_ack_1, ack => convTransposeD_CP_8453_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_update_start_
      -- CP-element group 22: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_Update/cr
      -- 
    ra_8642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3338_inst_ack_0, ack => convTransposeD_CP_8453_elements(22)); -- 
    cr_8646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(22), ack => RPIPE_Block3_start_3338_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3338_Update/$exit
      -- 
    ca_8647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3338_inst_ack_1, ack => convTransposeD_CP_8453_elements(23)); -- 
    rr_8655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(23), ack => type_cast_3342_inst_req_0); -- 
    rr_8669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(23), ack => RPIPE_Block3_start_3350_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_sample_completed_
      -- 
    ra_8656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3342_inst_ack_0, ack => convTransposeD_CP_8453_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	102 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3342_update_completed_
      -- 
    ca_8661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3342_inst_ack_1, ack => convTransposeD_CP_8453_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_update_start_
      -- CP-element group 26: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_sample_completed_
      -- 
    ra_8670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3350_inst_ack_0, ack => convTransposeD_CP_8453_elements(26)); -- 
    cr_8674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(26), ack => RPIPE_Block3_start_3350_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3350_Update/ca
      -- 
    ca_8675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3350_inst_ack_1, ack => convTransposeD_CP_8453_elements(27)); -- 
    rr_8683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(27), ack => RPIPE_Block3_start_3353_inst_req_0); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_update_start_
      -- 
    ra_8684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3353_inst_ack_0, ack => convTransposeD_CP_8453_elements(28)); -- 
    cr_8688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(28), ack => RPIPE_Block3_start_3353_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3353_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_Sample/rr
      -- 
    ca_8689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3353_inst_ack_1, ack => convTransposeD_CP_8453_elements(29)); -- 
    rr_8697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(29), ack => RPIPE_Block3_start_3356_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_update_start_
      -- CP-element group 30: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_Update/cr
      -- 
    ra_8698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3356_inst_ack_0, ack => convTransposeD_CP_8453_elements(30)); -- 
    cr_8702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(30), ack => RPIPE_Block3_start_3356_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3356_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_Sample/rr
      -- 
    ca_8703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3356_inst_ack_1, ack => convTransposeD_CP_8453_elements(31)); -- 
    rr_8725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(31), ack => RPIPE_Block3_start_3369_inst_req_0); -- 
    rr_8711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(31), ack => type_cast_3360_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_Sample/ra
      -- 
    ra_8712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3360_inst_ack_0, ack => convTransposeD_CP_8453_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	102 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3360_Update/ca
      -- 
    ca_8717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3360_inst_ack_1, ack => convTransposeD_CP_8453_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_update_start_
      -- CP-element group 34: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_Update/cr
      -- 
    ra_8726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3369_inst_ack_0, ack => convTransposeD_CP_8453_elements(34)); -- 
    cr_8730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(34), ack => RPIPE_Block3_start_3369_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3369_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_Sample/rr
      -- 
    ca_8731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3369_inst_ack_1, ack => convTransposeD_CP_8453_elements(35)); -- 
    rr_8739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(35), ack => type_cast_3373_inst_req_0); -- 
    rr_8753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(35), ack => RPIPE_Block3_start_3381_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_Sample/ra
      -- 
    ra_8740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3373_inst_ack_0, ack => convTransposeD_CP_8453_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	102 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3373_Update/ca
      -- 
    ca_8745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3373_inst_ack_1, ack => convTransposeD_CP_8453_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_update_start_
      -- CP-element group 38: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_Update/cr
      -- 
    ra_8754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3381_inst_ack_0, ack => convTransposeD_CP_8453_elements(38)); -- 
    cr_8758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(38), ack => RPIPE_Block3_start_3381_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	42 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3381_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_Sample/rr
      -- 
    ca_8759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3381_inst_ack_1, ack => convTransposeD_CP_8453_elements(39)); -- 
    rr_8781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(39), ack => RPIPE_Block3_start_3394_inst_req_0); -- 
    rr_8767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(39), ack => type_cast_3385_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_Sample/ra
      -- 
    ra_8768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3385_inst_ack_0, ack => convTransposeD_CP_8453_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	102 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3385_Update/ca
      -- 
    ca_8773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3385_inst_ack_1, ack => convTransposeD_CP_8453_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_update_start_
      -- CP-element group 42: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_Update/cr
      -- 
    ra_8782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3394_inst_ack_0, ack => convTransposeD_CP_8453_elements(42)); -- 
    cr_8786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(42), ack => RPIPE_Block3_start_3394_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	46 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3394_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_Sample/rr
      -- 
    ca_8787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3394_inst_ack_1, ack => convTransposeD_CP_8453_elements(43)); -- 
    rr_8809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(43), ack => RPIPE_Block3_start_3406_inst_req_0); -- 
    rr_8795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(43), ack => type_cast_3398_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_Sample/ra
      -- 
    ra_8796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3398_inst_ack_0, ack => convTransposeD_CP_8453_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	102 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3398_Update/ca
      -- 
    ca_8801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3398_inst_ack_1, ack => convTransposeD_CP_8453_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_update_start_
      -- CP-element group 46: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_Update/cr
      -- 
    ra_8810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3406_inst_ack_0, ack => convTransposeD_CP_8453_elements(46)); -- 
    cr_8814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(46), ack => RPIPE_Block3_start_3406_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3406_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_Sample/rr
      -- 
    ca_8815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3406_inst_ack_1, ack => convTransposeD_CP_8453_elements(47)); -- 
    rr_8823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(47), ack => RPIPE_Block3_start_3409_inst_req_0); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_update_start_
      -- CP-element group 48: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_Update/cr
      -- 
    ra_8824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3409_inst_ack_0, ack => convTransposeD_CP_8453_elements(48)); -- 
    cr_8828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(48), ack => RPIPE_Block3_start_3409_inst_req_1); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3409_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_Sample/rr
      -- 
    ca_8829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3409_inst_ack_1, ack => convTransposeD_CP_8453_elements(49)); -- 
    rr_8837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(49), ack => RPIPE_Block3_start_3412_inst_req_0); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_update_start_
      -- CP-element group 50: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_Update/cr
      -- 
    ra_8838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3412_inst_ack_0, ack => convTransposeD_CP_8453_elements(50)); -- 
    cr_8842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(50), ack => RPIPE_Block3_start_3412_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3412_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_Sample/rr
      -- 
    ca_8843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3412_inst_ack_1, ack => convTransposeD_CP_8453_elements(51)); -- 
    rr_8865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(51), ack => RPIPE_Block3_start_3425_inst_req_0); -- 
    rr_8851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(51), ack => type_cast_3416_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_Sample/ra
      -- 
    ra_8852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3416_inst_ack_0, ack => convTransposeD_CP_8453_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	0 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	102 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3416_Update/ca
      -- 
    ca_8857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3416_inst_ack_1, ack => convTransposeD_CP_8453_elements(53)); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	51 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_update_start_
      -- CP-element group 54: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_Update/cr
      -- 
    ra_8866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3425_inst_ack_0, ack => convTransposeD_CP_8453_elements(54)); -- 
    cr_8870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(54), ack => RPIPE_Block3_start_3425_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3425_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_Sample/rr
      -- 
    ca_8871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3425_inst_ack_1, ack => convTransposeD_CP_8453_elements(55)); -- 
    rr_8893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(55), ack => RPIPE_Block3_start_3437_inst_req_0); -- 
    rr_8879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(55), ack => type_cast_3429_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_Sample/ra
      -- 
    ra_8880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3429_inst_ack_0, ack => convTransposeD_CP_8453_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	0 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	102 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3429_Update/ca
      -- 
    ca_8885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3429_inst_ack_1, ack => convTransposeD_CP_8453_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_update_start_
      -- CP-element group 58: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_Update/cr
      -- 
    ra_8894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3437_inst_ack_0, ack => convTransposeD_CP_8453_elements(58)); -- 
    cr_8898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(58), ack => RPIPE_Block3_start_3437_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (9) 
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3437_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_Sample/rr
      -- 
    ca_8899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3437_inst_ack_1, ack => convTransposeD_CP_8453_elements(59)); -- 
    rr_8921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(59), ack => RPIPE_Block3_start_3450_inst_req_0); -- 
    rr_8907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(59), ack => type_cast_3441_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_Sample/ra
      -- 
    ra_8908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3441_inst_ack_0, ack => convTransposeD_CP_8453_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	0 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	102 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3441_Update/ca
      -- 
    ca_8913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3441_inst_ack_1, ack => convTransposeD_CP_8453_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_update_start_
      -- CP-element group 62: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_Update/cr
      -- 
    ra_8922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3450_inst_ack_0, ack => convTransposeD_CP_8453_elements(62)); -- 
    cr_8926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(62), ack => RPIPE_Block3_start_3450_inst_req_1); -- 
    -- CP-element group 63:  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3450_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_Sample/rr
      -- 
    ca_8927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3450_inst_ack_1, ack => convTransposeD_CP_8453_elements(63)); -- 
    rr_8949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(63), ack => RPIPE_Block3_start_3462_inst_req_0); -- 
    rr_8935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(63), ack => type_cast_3454_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_Sample/ra
      -- 
    ra_8936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3454_inst_ack_0, ack => convTransposeD_CP_8453_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	102 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3454_Update/ca
      -- 
    ca_8941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3454_inst_ack_1, ack => convTransposeD_CP_8453_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_update_start_
      -- CP-element group 66: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_Update/cr
      -- 
    ra_8950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3462_inst_ack_0, ack => convTransposeD_CP_8453_elements(66)); -- 
    cr_8954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(66), ack => RPIPE_Block3_start_3462_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	70 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3462_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_Sample/rr
      -- 
    ca_8955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3462_inst_ack_1, ack => convTransposeD_CP_8453_elements(67)); -- 
    rr_8977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(67), ack => RPIPE_Block3_start_3475_inst_req_0); -- 
    rr_8963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(67), ack => type_cast_3466_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_Sample/ra
      -- 
    ra_8964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3466_inst_ack_0, ack => convTransposeD_CP_8453_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	102 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3466_Update/ca
      -- 
    ca_8969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3466_inst_ack_1, ack => convTransposeD_CP_8453_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_update_start_
      -- CP-element group 70: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_Update/cr
      -- 
    ra_8978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3475_inst_ack_0, ack => convTransposeD_CP_8453_elements(70)); -- 
    cr_8982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(70), ack => RPIPE_Block3_start_3475_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	74 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3475_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_Sample/rr
      -- 
    ca_8983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3475_inst_ack_1, ack => convTransposeD_CP_8453_elements(71)); -- 
    rr_9005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(71), ack => RPIPE_Block3_start_3493_inst_req_0); -- 
    rr_8991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(71), ack => type_cast_3479_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_Sample/ra
      -- 
    ra_8992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3479_inst_ack_0, ack => convTransposeD_CP_8453_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	102 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3479_Update/ca
      -- 
    ca_8997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3479_inst_ack_1, ack => convTransposeD_CP_8453_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	71 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_update_start_
      -- CP-element group 74: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_Update/cr
      -- 
    ra_9006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3493_inst_ack_0, ack => convTransposeD_CP_8453_elements(74)); -- 
    cr_9010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(74), ack => RPIPE_Block3_start_3493_inst_req_1); -- 
    -- CP-element group 75:  fork  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (9) 
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3493_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_Sample/rr
      -- 
    ca_9011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3493_inst_ack_1, ack => convTransposeD_CP_8453_elements(75)); -- 
    rr_9033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(75), ack => RPIPE_Block3_start_3511_inst_req_0); -- 
    rr_9019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(75), ack => type_cast_3497_inst_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_Sample/ra
      -- 
    ra_9020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3497_inst_ack_0, ack => convTransposeD_CP_8453_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	102 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3497_Update/ca
      -- 
    ca_9025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3497_inst_ack_1, ack => convTransposeD_CP_8453_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_update_start_
      -- CP-element group 78: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_Update/cr
      -- 
    ra_9034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3511_inst_ack_0, ack => convTransposeD_CP_8453_elements(78)); -- 
    cr_9038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(78), ack => RPIPE_Block3_start_3511_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3511_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_Sample/rr
      -- 
    ca_9039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3511_inst_ack_1, ack => convTransposeD_CP_8453_elements(79)); -- 
    rr_9061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(79), ack => RPIPE_Block3_start_3523_inst_req_0); -- 
    rr_9047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(79), ack => type_cast_3515_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_Sample/ra
      -- 
    ra_9048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3515_inst_ack_0, ack => convTransposeD_CP_8453_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	102 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3515_Update/ca
      -- 
    ca_9053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3515_inst_ack_1, ack => convTransposeD_CP_8453_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_update_start_
      -- CP-element group 82: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_Update/cr
      -- 
    ra_9062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3523_inst_ack_0, ack => convTransposeD_CP_8453_elements(82)); -- 
    cr_9066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(82), ack => RPIPE_Block3_start_3523_inst_req_1); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3523_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_Sample/rr
      -- 
    ca_9067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3523_inst_ack_1, ack => convTransposeD_CP_8453_elements(83)); -- 
    rr_9075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(83), ack => RPIPE_Block3_start_3526_inst_req_0); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_update_start_
      -- CP-element group 84: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_Update/cr
      -- 
    ra_9076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3526_inst_ack_0, ack => convTransposeD_CP_8453_elements(84)); -- 
    cr_9080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(84), ack => RPIPE_Block3_start_3526_inst_req_1); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3526_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_Sample/rr
      -- 
    ca_9081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3526_inst_ack_1, ack => convTransposeD_CP_8453_elements(85)); -- 
    rr_9089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(85), ack => RPIPE_Block3_start_3529_inst_req_0); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_update_start_
      -- CP-element group 86: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_Sample/ra
      -- 
    ra_9090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3529_inst_ack_0, ack => convTransposeD_CP_8453_elements(86)); -- 
    cr_9094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(86), ack => RPIPE_Block3_start_3529_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3529_update_completed_
      -- 
    ca_9095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3529_inst_ack_1, ack => convTransposeD_CP_8453_elements(87)); -- 
    rr_9103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(87), ack => type_cast_3533_inst_req_0); -- 
    rr_9117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(87), ack => RPIPE_Block3_start_3542_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_Sample/$exit
      -- 
    ra_9104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3533_inst_ack_0, ack => convTransposeD_CP_8453_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	102 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3533_update_completed_
      -- 
    ca_9109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3533_inst_ack_1, ack => convTransposeD_CP_8453_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_update_start_
      -- CP-element group 90: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_Update/cr
      -- CP-element group 90: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_Sample/$exit
      -- 
    ra_9118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3542_inst_ack_0, ack => convTransposeD_CP_8453_elements(90)); -- 
    cr_9122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(90), ack => RPIPE_Block3_start_3542_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3542_Update/$exit
      -- 
    ca_9123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3542_inst_ack_1, ack => convTransposeD_CP_8453_elements(91)); -- 
    rr_9131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(91), ack => type_cast_3546_inst_req_0); -- 
    rr_9145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(91), ack => RPIPE_Block3_start_3554_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_sample_completed_
      -- 
    ra_9132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3546_inst_ack_0, ack => convTransposeD_CP_8453_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	102 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3546_update_completed_
      -- 
    ca_9137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3546_inst_ack_1, ack => convTransposeD_CP_8453_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_update_start_
      -- CP-element group 94: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_Sample/ra
      -- 
    ra_9146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3554_inst_ack_0, ack => convTransposeD_CP_8453_elements(94)); -- 
    cr_9150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(94), ack => RPIPE_Block3_start_3554_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3554_Update/$exit
      -- 
    ca_9151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3554_inst_ack_1, ack => convTransposeD_CP_8453_elements(95)); -- 
    rr_9159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(95), ack => type_cast_3558_inst_req_0); -- 
    rr_9173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(95), ack => RPIPE_Block3_start_3567_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_sample_completed_
      -- 
    ra_9160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3558_inst_ack_0, ack => convTransposeD_CP_8453_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	102 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3558_update_completed_
      -- 
    ca_9165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3558_inst_ack_1, ack => convTransposeD_CP_8453_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_update_start_
      -- CP-element group 98: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_sample_completed_
      -- 
    ra_9174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3567_inst_ack_0, ack => convTransposeD_CP_8453_elements(98)); -- 
    cr_9178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(98), ack => RPIPE_Block3_start_3567_inst_req_1); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/RPIPE_Block3_start_3567_update_completed_
      -- 
    ca_9179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_3567_inst_ack_1, ack => convTransposeD_CP_8453_elements(99)); -- 
    rr_9187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(99), ack => type_cast_3571_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_sample_completed_
      -- 
    ra_9188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3571_inst_ack_0, ack => convTransposeD_CP_8453_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/type_cast_3571_update_completed_
      -- 
    ca_9193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3571_inst_ack_1, ack => convTransposeD_CP_8453_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	81 
    -- CP-element group 102: 	69 
    -- CP-element group 102: 	77 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	97 
    -- CP-element group 102: 	61 
    -- CP-element group 102: 	93 
    -- CP-element group 102: 	101 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	41 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	37 
    -- CP-element group 102: 	33 
    -- CP-element group 102: 	73 
    -- CP-element group 102: 	89 
    -- CP-element group 102: 	5 
    -- CP-element group 102: 	9 
    -- CP-element group 102: 	13 
    -- CP-element group 102: 	17 
    -- CP-element group 102: 	21 
    -- CP-element group 102: 	25 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	138 
    -- CP-element group 102: 	139 
    -- CP-element group 102: 	142 
    -- CP-element group 102: 	141 
    -- CP-element group 102: 	143 
    -- CP-element group 102:  members (22) 
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody
      -- CP-element group 102: 	 branch_block_stmt_3273/assign_stmt_3584_to_assign_stmt_3617__exit__
      -- CP-element group 102: 	 branch_block_stmt_3273/assign_stmt_3584_to_assign_stmt_3617__entry__
      -- CP-element group 102: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577__exit__
      -- CP-element group 102: 	 branch_block_stmt_3273/assign_stmt_3276_to_assign_stmt_3577/$exit
      -- CP-element group 102: 	 branch_block_stmt_3273/assign_stmt_3584_to_assign_stmt_3617/$exit
      -- CP-element group 102: 	 branch_block_stmt_3273/assign_stmt_3584_to_assign_stmt_3617/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/Update/cr
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3634/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3627/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3620/$entry
      -- CP-element group 102: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/$entry
      -- 
    rr_9572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(102), ack => type_cast_3646_inst_req_0); -- 
    cr_9577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(102), ack => type_cast_3646_inst_req_1); -- 
    convTransposeD_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(81) & convTransposeD_CP_8453_elements(69) & convTransposeD_CP_8453_elements(77) & convTransposeD_CP_8453_elements(65) & convTransposeD_CP_8453_elements(57) & convTransposeD_CP_8453_elements(97) & convTransposeD_CP_8453_elements(61) & convTransposeD_CP_8453_elements(93) & convTransposeD_CP_8453_elements(101) & convTransposeD_CP_8453_elements(53) & convTransposeD_CP_8453_elements(41) & convTransposeD_CP_8453_elements(45) & convTransposeD_CP_8453_elements(37) & convTransposeD_CP_8453_elements(33) & convTransposeD_CP_8453_elements(73) & convTransposeD_CP_8453_elements(89) & convTransposeD_CP_8453_elements(5) & convTransposeD_CP_8453_elements(9) & convTransposeD_CP_8453_elements(13) & convTransposeD_CP_8453_elements(17) & convTransposeD_CP_8453_elements(21) & convTransposeD_CP_8453_elements(25);
      gj_convTransposeD_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	163 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_sample_completed_
      -- 
    ra_9208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3681_inst_ack_0, ack => convTransposeD_CP_8453_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	163 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	117 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_update_completed_
      -- 
    ca_9213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3681_inst_ack_1, ack => convTransposeD_CP_8453_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	163 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_Sample/ra
      -- 
    ra_9222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3685_inst_ack_0, ack => convTransposeD_CP_8453_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	163 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	117 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_Update/$exit
      -- 
    ca_9227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3685_inst_ack_1, ack => convTransposeD_CP_8453_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	163 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_sample_completed_
      -- 
    ra_9236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3689_inst_ack_0, ack => convTransposeD_CP_8453_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	163 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	117 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_update_completed_
      -- 
    ca_9241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3689_inst_ack_1, ack => convTransposeD_CP_8453_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	163 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_sample_completed_
      -- 
    ra_9250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3719_inst_ack_0, ack => convTransposeD_CP_8453_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	163 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (16) 
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_scale_1/$exit
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_scale_1/$entry
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_scale_1/scale_rename_ack
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_resize_1/$entry
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_resize_1/index_resize_ack
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_resize_1/$exit
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_scale_1/scale_rename_req
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_resize_1/index_resize_req
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_computed_1
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_scaled_1
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_index_resized_1
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_Sample/req
      -- 
    ca_9255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3719_inst_ack_1, ack => convTransposeD_CP_8453_elements(110)); -- 
    req_9280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(110), ack => array_obj_ref_3725_index_offset_req_0); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	127 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_sample_complete
      -- CP-element group 111: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_Sample/ack
      -- CP-element group 111: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_Sample/$exit
      -- 
    ack_9281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3725_index_offset_ack_0, ack => convTransposeD_CP_8453_elements(111)); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	163 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (11) 
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_offset_calculated
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_root_address_calculated
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_request/req
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_request/$entry
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_base_plus_offset/sum_rename_ack
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_base_plus_offset/sum_rename_req
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_base_plus_offset/$exit
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_base_plus_offset/$entry
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_Update/ack
      -- CP-element group 112: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_Update/$exit
      -- 
    ack_9286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3725_index_offset_ack_1, ack => convTransposeD_CP_8453_elements(112)); -- 
    req_9295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(112), ack => addr_of_3726_final_reg_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_request/ack
      -- CP-element group 113: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_request/$exit
      -- 
    ack_9296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3726_final_reg_ack_0, ack => convTransposeD_CP_8453_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	163 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (24) 
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Sample/word_access_start/word_0/$entry
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_plus_offset/sum_rename_ack
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_plus_offset/$entry
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_plus_offset/sum_rename_req
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Sample/word_access_start/word_0/rr
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_address_resized
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_word_addrgen/$exit
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_plus_offset/$exit
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_word_addrgen/$entry
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_addr_resize/base_resize_req
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_addr_resize/$entry
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_addr_resize/base_resize_ack
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_word_addrgen/root_register_req
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Sample/word_access_start/$entry
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_addr_resize/$exit
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_word_addrgen/root_register_ack
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_root_address_calculated
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_word_address_calculated
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_base_address_calculated
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_complete/ack
      -- CP-element group 114: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_complete/$exit
      -- 
    ack_9301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3726_final_reg_ack_1, ack => convTransposeD_CP_8453_elements(114)); -- 
    rr_9334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(114), ack => ptr_deref_3730_load_0_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Sample/word_access_start/word_0/ra
      -- CP-element group 115: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Sample/word_access_start/word_0/$exit
      -- CP-element group 115: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Sample/word_access_start/$exit
      -- CP-element group 115: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_sample_completed_
      -- 
    ra_9335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3730_load_0_ack_0, ack => convTransposeD_CP_8453_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	163 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	122 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/ptr_deref_3730_Merge/merge_ack
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/ptr_deref_3730_Merge/merge_req
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/ptr_deref_3730_Merge/$exit
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/ptr_deref_3730_Merge/$entry
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/word_access_complete/word_0/ca
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/word_access_complete/word_0/$exit
      -- CP-element group 116: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/word_access_complete/$exit
      -- 
    ca_9346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3730_load_0_ack_1, ack => convTransposeD_CP_8453_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	104 
    -- CP-element group 117: 	108 
    -- CP-element group 117: 	106 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (13) 
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_scale_1/$entry
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_Sample/req
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_scale_1/scale_rename_ack
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_scale_1/scale_rename_req
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_scale_1/$exit
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_resize_1/index_resize_ack
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_resize_1/index_resize_req
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_resize_1/$exit
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_resize_1/$entry
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_computed_1
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_scaled_1
      -- CP-element group 117: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_index_resized_1
      -- 
    req_9376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(117), ack => array_obj_ref_3748_index_offset_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(104) & convTransposeD_CP_8453_elements(108) & convTransposeD_CP_8453_elements(106);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	127 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_Sample/ack
      -- CP-element group 118: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_sample_complete
      -- 
    ack_9377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3748_index_offset_ack_0, ack => convTransposeD_CP_8453_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	163 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (11) 
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_offset_calculated
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_root_address_calculated
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_request/req
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_request/$entry
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_base_plus_offset/sum_rename_ack
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_base_plus_offset/sum_rename_req
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_base_plus_offset/$exit
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_base_plus_offset/$entry
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_Update/ack
      -- CP-element group 119: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_Update/$exit
      -- 
    ack_9382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3748_index_offset_ack_1, ack => convTransposeD_CP_8453_elements(119)); -- 
    req_9391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(119), ack => addr_of_3749_final_reg_req_0); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_request/ack
      -- CP-element group 120: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_request/$exit
      -- CP-element group 120: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_sample_completed_
      -- 
    ack_9392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3749_final_reg_ack_0, ack => convTransposeD_CP_8453_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	163 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (19) 
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_word_addrgen/$entry
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_word_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_word_addrgen/$exit
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_word_addrgen/root_register_req
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_plus_offset/$exit
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_plus_offset/sum_rename_req
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_complete/$exit
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_plus_offset/sum_rename_ack
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_complete/ack
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_root_address_calculated
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_plus_offset/$entry
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_addr_resize/base_resize_ack
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_addr_resize/base_resize_req
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_addr_resize/$exit
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_word_addrgen/root_register_ack
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_addr_resize/$entry
      -- CP-element group 121: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_base_address_resized
      -- 
    ack_9397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3749_final_reg_ack_1, ack => convTransposeD_CP_8453_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: 	116 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (9) 
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/word_access_start/word_0/$entry
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/word_access_start/word_0/rr
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/ptr_deref_3752_Split/$entry
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/word_access_start/$entry
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/ptr_deref_3752_Split/split_ack
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/ptr_deref_3752_Split/split_req
      -- CP-element group 122: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/ptr_deref_3752_Split/$exit
      -- 
    rr_9435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(122), ack => ptr_deref_3752_store_0_req_0); -- 
    convTransposeD_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(121) & convTransposeD_CP_8453_elements(116);
      gj_convTransposeD_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (5) 
      -- CP-element group 123: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/word_access_start/word_0/$exit
      -- CP-element group 123: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/word_access_start/word_0/ra
      -- CP-element group 123: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/word_access_start/$exit
      -- CP-element group 123: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Sample/$exit
      -- 
    ra_9436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3752_store_0_ack_0, ack => convTransposeD_CP_8453_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	163 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Update/word_access_complete/$exit
      -- CP-element group 124: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Update/word_access_complete/word_0/ca
      -- CP-element group 124: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Update/word_access_complete/word_0/$exit
      -- 
    ca_9447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3752_store_0_ack_1, ack => convTransposeD_CP_8453_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	163 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_Sample/ra
      -- 
    ra_9456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3757_inst_ack_0, ack => convTransposeD_CP_8453_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	163 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_Update/ca
      -- 
    ca_9461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3757_inst_ack_1, ack => convTransposeD_CP_8453_elements(126)); -- 
    -- CP-element group 127:  branch  join  transition  place  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	111 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	118 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (10) 
      -- CP-element group 127: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769__exit__
      -- CP-element group 127: 	 branch_block_stmt_3273/if_stmt_3770__entry__
      -- CP-element group 127: 	 branch_block_stmt_3273/R_cmp_3771_place
      -- CP-element group 127: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/$exit
      -- CP-element group 127: 	 branch_block_stmt_3273/if_stmt_3770_dead_link/$entry
      -- CP-element group 127: 	 branch_block_stmt_3273/if_stmt_3770_eval_test/$entry
      -- CP-element group 127: 	 branch_block_stmt_3273/if_stmt_3770_eval_test/$exit
      -- CP-element group 127: 	 branch_block_stmt_3273/if_stmt_3770_eval_test/branch_req
      -- CP-element group 127: 	 branch_block_stmt_3273/if_stmt_3770_if_link/$entry
      -- CP-element group 127: 	 branch_block_stmt_3273/if_stmt_3770_else_link/$entry
      -- 
    branch_req_9469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(127), ack => if_stmt_3770_branch_req_0); -- 
    convTransposeD_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(111) & convTransposeD_CP_8453_elements(124) & convTransposeD_CP_8453_elements(118) & convTransposeD_CP_8453_elements(126);
      gj_convTransposeD_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	178 
    -- CP-element group 128: 	179 
    -- CP-element group 128: 	172 
    -- CP-element group 128: 	173 
    -- CP-element group 128: 	175 
    -- CP-element group 128: 	176 
    -- CP-element group 128:  members (40) 
      -- CP-element group 128: 	 branch_block_stmt_3273/assign_stmt_3782__exit__
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258
      -- CP-element group 128: 	 branch_block_stmt_3273/assign_stmt_3782__entry__
      -- CP-element group 128: 	 branch_block_stmt_3273/merge_stmt_3776__exit__
      -- CP-element group 128: 	 branch_block_stmt_3273/whilex_xbody_ifx_xthen
      -- CP-element group 128: 	 branch_block_stmt_3273/if_stmt_3770_if_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_3273/if_stmt_3770_if_link/if_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_3273/assign_stmt_3782/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/assign_stmt_3782/$exit
      -- CP-element group 128: 	 branch_block_stmt_3273/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 128: 	 branch_block_stmt_3273/merge_stmt_3776_PhiReqMerge
      -- CP-element group 128: 	 branch_block_stmt_3273/merge_stmt_3776_PhiAck/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/merge_stmt_3776_PhiAck/$exit
      -- CP-element group 128: 	 branch_block_stmt_3273/merge_stmt_3776_PhiAck/dummy
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/Update/cr
      -- 
    if_choice_transition_9474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3770_branch_ack_1, ack => convTransposeD_CP_8453_elements(128)); -- 
    rr_9806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(128), ack => type_cast_3844_inst_req_0); -- 
    cr_9811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(128), ack => type_cast_3844_inst_req_1); -- 
    rr_9829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(128), ack => type_cast_3838_inst_req_0); -- 
    cr_9834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(128), ack => type_cast_3838_inst_req_1); -- 
    rr_9852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(128), ack => type_cast_3834_inst_req_0); -- 
    cr_9857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(128), ack => type_cast_3834_inst_req_1); -- 
    -- CP-element group 129:  fork  transition  place  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	133 
    -- CP-element group 129: 	130 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (21) 
      -- CP-element group 129: 	 branch_block_stmt_3273/merge_stmt_3784__exit__
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820__entry__
      -- CP-element group 129: 	 branch_block_stmt_3273/whilex_xbody_ifx_xelse
      -- CP-element group 129: 	 branch_block_stmt_3273/if_stmt_3770_else_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_3273/if_stmt_3770_else_link/else_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/$entry
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_update_start_
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_Sample/rr
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_update_start_
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_Update/cr
      -- CP-element group 129: 	 branch_block_stmt_3273/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_3273/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 129: 	 branch_block_stmt_3273/merge_stmt_3784_PhiReqMerge
      -- CP-element group 129: 	 branch_block_stmt_3273/merge_stmt_3784_PhiAck/$entry
      -- CP-element group 129: 	 branch_block_stmt_3273/merge_stmt_3784_PhiAck/$exit
      -- CP-element group 129: 	 branch_block_stmt_3273/merge_stmt_3784_PhiAck/dummy
      -- 
    else_choice_transition_9478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3770_branch_ack_0, ack => convTransposeD_CP_8453_elements(129)); -- 
    rr_9494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(129), ack => type_cast_3793_inst_req_0); -- 
    cr_9499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(129), ack => type_cast_3793_inst_req_1); -- 
    cr_9513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(129), ack => type_cast_3802_inst_req_1); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_Sample/ra
      -- 
    ra_9495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3793_inst_ack_0, ack => convTransposeD_CP_8453_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3793_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_Sample/rr
      -- 
    ca_9500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3793_inst_ack_1, ack => convTransposeD_CP_8453_elements(131)); -- 
    rr_9508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(131), ack => type_cast_3802_inst_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_Sample/ra
      -- 
    ra_9509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3802_inst_ack_0, ack => convTransposeD_CP_8453_elements(132)); -- 
    -- CP-element group 133:  branch  transition  place  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	129 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (13) 
      -- CP-element group 133: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820__exit__
      -- CP-element group 133: 	 branch_block_stmt_3273/if_stmt_3821__entry__
      -- CP-element group 133: 	 branch_block_stmt_3273/R_cmp247_3822_place
      -- CP-element group 133: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/$exit
      -- CP-element group 133: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_3273/assign_stmt_3790_to_assign_stmt_3820/type_cast_3802_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_3273/if_stmt_3821_dead_link/$entry
      -- CP-element group 133: 	 branch_block_stmt_3273/if_stmt_3821_eval_test/$entry
      -- CP-element group 133: 	 branch_block_stmt_3273/if_stmt_3821_eval_test/$exit
      -- CP-element group 133: 	 branch_block_stmt_3273/if_stmt_3821_eval_test/branch_req
      -- CP-element group 133: 	 branch_block_stmt_3273/if_stmt_3821_if_link/$entry
      -- CP-element group 133: 	 branch_block_stmt_3273/if_stmt_3821_else_link/$entry
      -- 
    ca_9514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3802_inst_ack_1, ack => convTransposeD_CP_8453_elements(133)); -- 
    branch_req_9522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_9522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(133), ack => if_stmt_3821_branch_req_0); -- 
    -- CP-element group 134:  transition  place  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (15) 
      -- CP-element group 134: 	 branch_block_stmt_3273/merge_stmt_3855__exit__
      -- CP-element group 134: 	 branch_block_stmt_3273/assign_stmt_3860__entry__
      -- CP-element group 134: 	 branch_block_stmt_3273/ifx_xelse_whilex_xend
      -- CP-element group 134: 	 branch_block_stmt_3273/if_stmt_3821_if_link/$exit
      -- CP-element group 134: 	 branch_block_stmt_3273/if_stmt_3821_if_link/if_choice_transition
      -- CP-element group 134: 	 branch_block_stmt_3273/assign_stmt_3860/$entry
      -- CP-element group 134: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_Sample/req
      -- CP-element group 134: 	 branch_block_stmt_3273/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 134: 	 branch_block_stmt_3273/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 134: 	 branch_block_stmt_3273/merge_stmt_3855_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_3273/merge_stmt_3855_PhiAck/$entry
      -- CP-element group 134: 	 branch_block_stmt_3273/merge_stmt_3855_PhiAck/$exit
      -- CP-element group 134: 	 branch_block_stmt_3273/merge_stmt_3855_PhiAck/dummy
      -- 
    if_choice_transition_9527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3821_branch_ack_1, ack => convTransposeD_CP_8453_elements(134)); -- 
    req_9547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(134), ack => WPIPE_Block3_done_3857_inst_req_0); -- 
    -- CP-element group 135:  fork  transition  place  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	168 
    -- CP-element group 135: 	170 
    -- CP-element group 135: 	165 
    -- CP-element group 135: 	167 
    -- CP-element group 135: 	164 
    -- CP-element group 135:  members (22) 
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258
      -- CP-element group 135: 	 branch_block_stmt_3273/if_stmt_3821_else_link/$exit
      -- CP-element group 135: 	 branch_block_stmt_3273/if_stmt_3821_else_link/else_choice_transition
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/Sample/rr
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/Update/cr
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/Sample/rr
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/Update/cr
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3828/$entry
      -- CP-element group 135: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/$entry
      -- 
    else_choice_transition_9531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3821_branch_ack_0, ack => convTransposeD_CP_8453_elements(135)); -- 
    rr_9749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(135), ack => type_cast_3846_inst_req_0); -- 
    cr_9754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(135), ack => type_cast_3846_inst_req_1); -- 
    rr_9772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(135), ack => type_cast_3840_inst_req_0); -- 
    cr_9777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(135), ack => type_cast_3840_inst_req_1); -- 
    -- CP-element group 136:  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (6) 
      -- CP-element group 136: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_update_start_
      -- CP-element group 136: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_Sample/ack
      -- CP-element group 136: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_Update/req
      -- 
    ack_9548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3857_inst_ack_0, ack => convTransposeD_CP_8453_elements(136)); -- 
    req_9552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(136), ack => WPIPE_Block3_done_3857_inst_req_1); -- 
    -- CP-element group 137:  transition  place  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (16) 
      -- CP-element group 137: 	 branch_block_stmt_3273/branch_block_stmt_3273__exit__
      -- CP-element group 137: 	 $exit
      -- CP-element group 137: 	 branch_block_stmt_3273/$exit
      -- CP-element group 137: 	 branch_block_stmt_3273/assign_stmt_3860__exit__
      -- CP-element group 137: 	 branch_block_stmt_3273/return__
      -- CP-element group 137: 	 branch_block_stmt_3273/merge_stmt_3862__exit__
      -- CP-element group 137: 	 branch_block_stmt_3273/assign_stmt_3860/$exit
      -- CP-element group 137: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_3273/assign_stmt_3860/WPIPE_Block3_done_3857_Update/ack
      -- CP-element group 137: 	 branch_block_stmt_3273/return___PhiReq/$entry
      -- CP-element group 137: 	 branch_block_stmt_3273/return___PhiReq/$exit
      -- CP-element group 137: 	 branch_block_stmt_3273/merge_stmt_3862_PhiReqMerge
      -- CP-element group 137: 	 branch_block_stmt_3273/merge_stmt_3862_PhiAck/$entry
      -- CP-element group 137: 	 branch_block_stmt_3273/merge_stmt_3862_PhiAck/$exit
      -- CP-element group 137: 	 branch_block_stmt_3273/merge_stmt_3862_PhiAck/dummy
      -- 
    ack_9553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3857_inst_ack_1, ack => convTransposeD_CP_8453_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	102 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/Sample/ra
      -- 
    ra_9573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3646_inst_ack_0, ack => convTransposeD_CP_8453_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	102 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/Update/ca
      -- 
    ca_9578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3646_inst_ack_1, ack => convTransposeD_CP_8453_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	144 
    -- CP-element group 140:  members (5) 
      -- CP-element group 140: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/$exit
      -- CP-element group 140: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/$exit
      -- CP-element group 140: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/$exit
      -- CP-element group 140: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3646/SplitProtocol/$exit
      -- CP-element group 140: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_req
      -- 
    phi_stmt_3641_req_9579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3641_req_9579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(140), ack => phi_stmt_3641_req_1); -- 
    convTransposeD_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(138) & convTransposeD_CP_8453_elements(139);
      gj_convTransposeD_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  transition  output  delay-element  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	102 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	144 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3634/$exit
      -- CP-element group 141: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/$exit
      -- CP-element group 141: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3638_konst_delay_trans
      -- CP-element group 141: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_req
      -- 
    phi_stmt_3634_req_9587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3634_req_9587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(141), ack => phi_stmt_3634_req_0); -- 
    -- Element group convTransposeD_CP_8453_elements(141) is a control-delay.
    cp_element_141_delay: control_delay_element  generic map(name => " 141_delay", delay_value => 1)  port map(req => convTransposeD_CP_8453_elements(102), ack => convTransposeD_CP_8453_elements(141), clk => clk, reset =>reset);
    -- CP-element group 142:  transition  output  delay-element  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	102 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3627/$exit
      -- CP-element group 142: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/$exit
      -- CP-element group 142: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3631_konst_delay_trans
      -- CP-element group 142: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_req
      -- 
    phi_stmt_3627_req_9595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3627_req_9595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(142), ack => phi_stmt_3627_req_0); -- 
    -- Element group convTransposeD_CP_8453_elements(142) is a control-delay.
    cp_element_142_delay: control_delay_element  generic map(name => " 142_delay", delay_value => 1)  port map(req => convTransposeD_CP_8453_elements(102), ack => convTransposeD_CP_8453_elements(142), clk => clk, reset =>reset);
    -- CP-element group 143:  transition  output  delay-element  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	102 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3620/$exit
      -- CP-element group 143: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/$exit
      -- CP-element group 143: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3624_konst_delay_trans
      -- CP-element group 143: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_req
      -- 
    phi_stmt_3620_req_9603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3620_req_9603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(143), ack => phi_stmt_3620_req_0); -- 
    -- Element group convTransposeD_CP_8453_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => convTransposeD_CP_8453_elements(102), ack => convTransposeD_CP_8453_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  join  transition  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: 	140 
    -- CP-element group 144: 	141 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	158 
    -- CP-element group 144:  members (1) 
      -- CP-element group 144: 	 branch_block_stmt_3273/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(142) & convTransposeD_CP_8453_elements(140) & convTransposeD_CP_8453_elements(141) & convTransposeD_CP_8453_elements(143);
      gj_convTransposeD_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	1 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/Sample/ra
      -- 
    ra_9623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3644_inst_ack_0, ack => convTransposeD_CP_8453_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	1 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/Update/ca
      -- 
    ca_9628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3644_inst_ack_1, ack => convTransposeD_CP_8453_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	157 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/$exit
      -- CP-element group 147: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/$exit
      -- CP-element group 147: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/$exit
      -- CP-element group 147: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_sources/type_cast_3644/SplitProtocol/$exit
      -- CP-element group 147: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3641/phi_stmt_3641_req
      -- 
    phi_stmt_3641_req_9629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3641_req_9629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(147), ack => phi_stmt_3641_req_0); -- 
    convTransposeD_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(145) & convTransposeD_CP_8453_elements(146);
      gj_convTransposeD_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	1 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (2) 
      -- CP-element group 148: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/Sample/ra
      -- 
    ra_9646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3640_inst_ack_0, ack => convTransposeD_CP_8453_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	1 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (2) 
      -- CP-element group 149: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/Update/ca
      -- 
    ca_9651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3640_inst_ack_1, ack => convTransposeD_CP_8453_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	157 
    -- CP-element group 150:  members (5) 
      -- CP-element group 150: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/$exit
      -- CP-element group 150: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/$exit
      -- CP-element group 150: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/$exit
      -- CP-element group 150: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_sources/type_cast_3640/SplitProtocol/$exit
      -- CP-element group 150: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3634/phi_stmt_3634_req
      -- 
    phi_stmt_3634_req_9652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3634_req_9652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(150), ack => phi_stmt_3634_req_1); -- 
    convTransposeD_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(148) & convTransposeD_CP_8453_elements(149);
      gj_convTransposeD_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	1 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (2) 
      -- CP-element group 151: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/Sample/ra
      -- 
    ra_9669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3633_inst_ack_0, ack => convTransposeD_CP_8453_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	1 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (2) 
      -- CP-element group 152: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/Update/ca
      -- 
    ca_9674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3633_inst_ack_1, ack => convTransposeD_CP_8453_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	157 
    -- CP-element group 153:  members (5) 
      -- CP-element group 153: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/$exit
      -- CP-element group 153: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/$exit
      -- CP-element group 153: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/$exit
      -- CP-element group 153: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_sources/type_cast_3633/SplitProtocol/$exit
      -- CP-element group 153: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3627/phi_stmt_3627_req
      -- 
    phi_stmt_3627_req_9675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3627_req_9675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(153), ack => phi_stmt_3627_req_1); -- 
    convTransposeD_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(151) & convTransposeD_CP_8453_elements(152);
      gj_convTransposeD_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	1 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (2) 
      -- CP-element group 154: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/Sample/ra
      -- 
    ra_9692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3626_inst_ack_0, ack => convTransposeD_CP_8453_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	1 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (2) 
      -- CP-element group 155: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/Update/ca
      -- 
    ca_9697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3626_inst_ack_1, ack => convTransposeD_CP_8453_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/$exit
      -- CP-element group 156: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/$exit
      -- CP-element group 156: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/$exit
      -- CP-element group 156: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_sources/type_cast_3626/SplitProtocol/$exit
      -- CP-element group 156: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/phi_stmt_3620/phi_stmt_3620_req
      -- 
    phi_stmt_3620_req_9698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3620_req_9698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(156), ack => phi_stmt_3620_req_1); -- 
    convTransposeD_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(154) & convTransposeD_CP_8453_elements(155);
      gj_convTransposeD_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	147 
    -- CP-element group 157: 	156 
    -- CP-element group 157: 	153 
    -- CP-element group 157: 	150 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_3273/ifx_xend258_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(147) & convTransposeD_CP_8453_elements(156) & convTransposeD_CP_8453_elements(153) & convTransposeD_CP_8453_elements(150);
      gj_convTransposeD_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  merge  fork  transition  place  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: 	144 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	162 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	160 
    -- CP-element group 158: 	161 
    -- CP-element group 158:  members (2) 
      -- CP-element group 158: 	 branch_block_stmt_3273/merge_stmt_3619_PhiReqMerge
      -- CP-element group 158: 	 branch_block_stmt_3273/merge_stmt_3619_PhiAck/$entry
      -- 
    convTransposeD_CP_8453_elements(158) <= OrReduce(convTransposeD_CP_8453_elements(157) & convTransposeD_CP_8453_elements(144));
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	163 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_3273/merge_stmt_3619_PhiAck/phi_stmt_3620_ack
      -- 
    phi_stmt_3620_ack_9703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3620_ack_0, ack => convTransposeD_CP_8453_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	163 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_3273/merge_stmt_3619_PhiAck/phi_stmt_3627_ack
      -- 
    phi_stmt_3627_ack_9704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3627_ack_0, ack => convTransposeD_CP_8453_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	158 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_3273/merge_stmt_3619_PhiAck/phi_stmt_3634_ack
      -- 
    phi_stmt_3634_ack_9705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3634_ack_0, ack => convTransposeD_CP_8453_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	158 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_3273/merge_stmt_3619_PhiAck/phi_stmt_3641_ack
      -- 
    phi_stmt_3641_ack_9706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3641_ack_0, ack => convTransposeD_CP_8453_elements(162)); -- 
    -- CP-element group 163:  join  fork  transition  place  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: 	159 
    -- CP-element group 163: 	160 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	103 
    -- CP-element group 163: 	104 
    -- CP-element group 163: 	110 
    -- CP-element group 163: 	109 
    -- CP-element group 163: 	107 
    -- CP-element group 163: 	108 
    -- CP-element group 163: 	105 
    -- CP-element group 163: 	121 
    -- CP-element group 163: 	106 
    -- CP-element group 163: 	119 
    -- CP-element group 163: 	116 
    -- CP-element group 163: 	114 
    -- CP-element group 163: 	124 
    -- CP-element group 163: 	112 
    -- CP-element group 163: 	125 
    -- CP-element group 163: 	126 
    -- CP-element group 163:  members (56) 
      -- CP-element group 163: 	 branch_block_stmt_3273/merge_stmt_3619__exit__
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769__entry__
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/word_access_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_update_start
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_complete/req
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3681_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3749_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Update/word_access_complete/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Update/word_access_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_complete/req
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/addr_of_3726_complete/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3752_Update/word_access_complete/word_0/cr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_Update/req
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3719_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3748_final_index_sum_regn_update_start
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_Update/req
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/word_access_complete/word_0/cr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/array_obj_ref_3725_final_index_sum_regn_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3689_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/ptr_deref_3730_Update/word_access_complete/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3685_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3273/assign_stmt_3653_to_assign_stmt_3769/type_cast_3757_Update/cr
      -- CP-element group 163: 	 branch_block_stmt_3273/merge_stmt_3619_PhiAck/$exit
      -- 
    rr_9221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3685_inst_req_0); -- 
    cr_9212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3681_inst_req_1); -- 
    rr_9207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3681_inst_req_0); -- 
    req_9396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => addr_of_3749_final_reg_req_1); -- 
    cr_9254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3719_inst_req_1); -- 
    req_9300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => addr_of_3726_final_reg_req_1); -- 
    cr_9446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => ptr_deref_3752_store_0_req_1); -- 
    rr_9249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3719_inst_req_0); -- 
    req_9381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => array_obj_ref_3748_index_offset_req_1); -- 
    cr_9240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3689_inst_req_1); -- 
    rr_9235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3689_inst_req_0); -- 
    req_9285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => array_obj_ref_3725_index_offset_req_1); -- 
    cr_9345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => ptr_deref_3730_load_0_req_1); -- 
    cr_9226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3685_inst_req_1); -- 
    rr_9455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3757_inst_req_0); -- 
    cr_9460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(163), ack => type_cast_3757_inst_req_1); -- 
    convTransposeD_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(162) & convTransposeD_CP_8453_elements(159) & convTransposeD_CP_8453_elements(160) & convTransposeD_CP_8453_elements(161);
      gj_convTransposeD_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	135 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/Sample/ra
      -- 
    ra_9750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3846_inst_ack_0, ack => convTransposeD_CP_8453_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	135 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/Update/ca
      -- 
    ca_9755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3846_inst_ack_1, ack => convTransposeD_CP_8453_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	171 
    -- CP-element group 166:  members (5) 
      -- CP-element group 166: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/$exit
      -- CP-element group 166: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/$exit
      -- CP-element group 166: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/$exit
      -- CP-element group 166: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3846/SplitProtocol/$exit
      -- CP-element group 166: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_req
      -- 
    phi_stmt_3841_req_9756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3841_req_9756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(166), ack => phi_stmt_3841_req_1); -- 
    convTransposeD_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(165) & convTransposeD_CP_8453_elements(164);
      gj_convTransposeD_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	135 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/Sample/ra
      -- 
    ra_9773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3840_inst_ack_0, ack => convTransposeD_CP_8453_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	135 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (2) 
      -- CP-element group 168: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/Update/ca
      -- 
    ca_9778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3840_inst_ack_1, ack => convTransposeD_CP_8453_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (5) 
      -- CP-element group 169: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/$exit
      -- CP-element group 169: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/$exit
      -- CP-element group 169: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/$exit
      -- CP-element group 169: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3840/SplitProtocol/$exit
      -- CP-element group 169: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_req
      -- 
    phi_stmt_3835_req_9779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3835_req_9779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(169), ack => phi_stmt_3835_req_1); -- 
    convTransposeD_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(168) & convTransposeD_CP_8453_elements(167);
      gj_convTransposeD_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  transition  output  delay-element  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	135 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3828/$exit
      -- CP-element group 170: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/$exit
      -- CP-element group 170: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3832_konst_delay_trans
      -- CP-element group 170: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_req
      -- 
    phi_stmt_3828_req_9787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3828_req_9787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(170), ack => phi_stmt_3828_req_0); -- 
    -- Element group convTransposeD_CP_8453_elements(170) is a control-delay.
    cp_element_170_delay: control_delay_element  generic map(name => " 170_delay", delay_value => 1)  port map(req => convTransposeD_CP_8453_elements(135), ack => convTransposeD_CP_8453_elements(170), clk => clk, reset =>reset);
    -- CP-element group 171:  join  transition  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: 	170 
    -- CP-element group 171: 	166 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	182 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 branch_block_stmt_3273/ifx_xelse_ifx_xend258_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(169) & convTransposeD_CP_8453_elements(170) & convTransposeD_CP_8453_elements(166);
      gj_convTransposeD_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	128 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/Sample/ra
      -- 
    ra_9807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3844_inst_ack_0, ack => convTransposeD_CP_8453_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	128 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (2) 
      -- CP-element group 173: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/Update/ca
      -- 
    ca_9812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3844_inst_ack_1, ack => convTransposeD_CP_8453_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	181 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/$exit
      -- CP-element group 174: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/$exit
      -- CP-element group 174: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/$exit
      -- CP-element group 174: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_sources/type_cast_3844/SplitProtocol/$exit
      -- CP-element group 174: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3841/phi_stmt_3841_req
      -- 
    phi_stmt_3841_req_9813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3841_req_9813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(174), ack => phi_stmt_3841_req_0); -- 
    convTransposeD_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(172) & convTransposeD_CP_8453_elements(173);
      gj_convTransposeD_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	128 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (2) 
      -- CP-element group 175: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/Sample/ra
      -- 
    ra_9830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3838_inst_ack_0, ack => convTransposeD_CP_8453_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	128 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/Update/ca
      -- 
    ca_9835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3838_inst_ack_1, ack => convTransposeD_CP_8453_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	181 
    -- CP-element group 177:  members (5) 
      -- CP-element group 177: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/$exit
      -- CP-element group 177: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/$exit
      -- CP-element group 177: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/$exit
      -- CP-element group 177: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_sources/type_cast_3838/SplitProtocol/$exit
      -- CP-element group 177: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3835/phi_stmt_3835_req
      -- 
    phi_stmt_3835_req_9836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3835_req_9836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(177), ack => phi_stmt_3835_req_0); -- 
    convTransposeD_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(175) & convTransposeD_CP_8453_elements(176);
      gj_convTransposeD_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	128 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/Sample/ra
      -- 
    ra_9853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3834_inst_ack_0, ack => convTransposeD_CP_8453_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	128 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/Update/ca
      -- 
    ca_9858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3834_inst_ack_1, ack => convTransposeD_CP_8453_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (5) 
      -- CP-element group 180: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/$exit
      -- CP-element group 180: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/$exit
      -- CP-element group 180: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/$exit
      -- CP-element group 180: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_sources/type_cast_3834/SplitProtocol/$exit
      -- CP-element group 180: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/phi_stmt_3828/phi_stmt_3828_req
      -- 
    phi_stmt_3828_req_9859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3828_req_9859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_8453_elements(180), ack => phi_stmt_3828_req_1); -- 
    convTransposeD_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(178) & convTransposeD_CP_8453_elements(179);
      gj_convTransposeD_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	174 
    -- CP-element group 181: 	177 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_3273/ifx_xthen_ifx_xend258_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(174) & convTransposeD_CP_8453_elements(177) & convTransposeD_CP_8453_elements(180);
      gj_convTransposeD_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  merge  fork  transition  place  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	171 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	185 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_3273/merge_stmt_3827_PhiReqMerge
      -- CP-element group 182: 	 branch_block_stmt_3273/merge_stmt_3827_PhiAck/$entry
      -- 
    convTransposeD_CP_8453_elements(182) <= OrReduce(convTransposeD_CP_8453_elements(171) & convTransposeD_CP_8453_elements(181));
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	186 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_3273/merge_stmt_3827_PhiAck/phi_stmt_3828_ack
      -- 
    phi_stmt_3828_ack_9864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3828_ack_0, ack => convTransposeD_CP_8453_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_3273/merge_stmt_3827_PhiAck/phi_stmt_3835_ack
      -- 
    phi_stmt_3835_ack_9865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3835_ack_0, ack => convTransposeD_CP_8453_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_3273/merge_stmt_3827_PhiAck/phi_stmt_3841_ack
      -- 
    phi_stmt_3841_ack_9866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3841_ack_0, ack => convTransposeD_CP_8453_elements(185)); -- 
    -- CP-element group 186:  join  transition  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: 	185 
    -- CP-element group 186: 	183 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	1 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_3273/merge_stmt_3827_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_8453_elements(184) & convTransposeD_CP_8453_elements(185) & convTransposeD_CP_8453_elements(183);
      gj_convTransposeD_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_8453_elements(186), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom217_3747_resized : std_logic_vector(13 downto 0);
    signal R_idxprom217_3747_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3724_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3724_scaled : std_logic_vector(13 downto 0);
    signal add103_3485 : std_logic_vector(31 downto 0);
    signal add108_3503 : std_logic_vector(31 downto 0);
    signal add113_3521 : std_logic_vector(31 downto 0);
    signal add135_3552 : std_logic_vector(63 downto 0);
    signal add147_3577 : std_logic_vector(63 downto 0);
    signal add158_3595 : std_logic_vector(15 downto 0);
    signal add16_3323 : std_logic_vector(31 downto 0);
    signal add176_3601 : std_logic_vector(15 downto 0);
    signal add189_3612 : std_logic_vector(15 downto 0);
    signal add208_3700 : std_logic_vector(63 downto 0);
    signal add210_3710 : std_logic_vector(63 downto 0);
    signal add222_3764 : std_logic_vector(31 downto 0);
    signal add229_3782 : std_logic_vector(15 downto 0);
    signal add28_3348 : std_logic_vector(31 downto 0);
    signal add52_3379 : std_logic_vector(15 downto 0);
    signal add64_3404 : std_logic_vector(15 downto 0);
    signal add86_3435 : std_logic_vector(15 downto 0);
    signal add95_3460 : std_logic_vector(15 downto 0);
    signal add_3298 : std_logic_vector(15 downto 0);
    signal add_src_0x_x0_3658 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3725_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3725_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3748_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3748_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3748_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3748_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3748_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3748_root_address : std_logic_vector(13 downto 0);
    signal arrayidx213_3727 : std_logic_vector(31 downto 0);
    signal arrayidx218_3750 : std_logic_vector(31 downto 0);
    signal call101_3476 : std_logic_vector(7 downto 0);
    signal call106_3494 : std_logic_vector(7 downto 0);
    signal call111_3512 : std_logic_vector(7 downto 0);
    signal call114_3524 : std_logic_vector(7 downto 0);
    signal call121_3527 : std_logic_vector(7 downto 0);
    signal call126_3530 : std_logic_vector(7 downto 0);
    signal call133_3543 : std_logic_vector(7 downto 0);
    signal call138_3555 : std_logic_vector(7 downto 0);
    signal call145_3568 : std_logic_vector(7 downto 0);
    signal call14_3314 : std_logic_vector(7 downto 0);
    signal call19_3326 : std_logic_vector(7 downto 0);
    signal call26_3339 : std_logic_vector(7 downto 0);
    signal call31_3351 : std_logic_vector(7 downto 0);
    signal call38_3354 : std_logic_vector(7 downto 0);
    signal call3_3289 : std_logic_vector(7 downto 0);
    signal call43_3357 : std_logic_vector(7 downto 0);
    signal call50_3370 : std_logic_vector(7 downto 0);
    signal call55_3382 : std_logic_vector(7 downto 0);
    signal call62_3395 : std_logic_vector(7 downto 0);
    signal call67_3407 : std_logic_vector(7 downto 0);
    signal call74_3410 : std_logic_vector(7 downto 0);
    signal call79_3413 : std_logic_vector(7 downto 0);
    signal call7_3301 : std_logic_vector(7 downto 0);
    signal call84_3426 : std_logic_vector(7 downto 0);
    signal call88_3438 : std_logic_vector(7 downto 0);
    signal call93_3451 : std_logic_vector(7 downto 0);
    signal call97_3463 : std_logic_vector(7 downto 0);
    signal call_3276 : std_logic_vector(7 downto 0);
    signal cmp237_3799 : std_logic_vector(0 downto 0);
    signal cmp247_3820 : std_logic_vector(0 downto 0);
    signal cmp_3769 : std_logic_vector(0 downto 0);
    signal conv102_3480 : std_logic_vector(31 downto 0);
    signal conv107_3498 : std_logic_vector(31 downto 0);
    signal conv112_3516 : std_logic_vector(31 downto 0);
    signal conv12_3305 : std_logic_vector(31 downto 0);
    signal conv131_3534 : std_logic_vector(63 downto 0);
    signal conv134_3547 : std_logic_vector(63 downto 0);
    signal conv143_3559 : std_logic_vector(63 downto 0);
    signal conv146_3572 : std_logic_vector(63 downto 0);
    signal conv15_3318 : std_logic_vector(31 downto 0);
    signal conv196_3682 : std_logic_vector(63 downto 0);
    signal conv201_3686 : std_logic_vector(63 downto 0);
    signal conv206_3690 : std_logic_vector(63 downto 0);
    signal conv221_3758 : std_logic_vector(31 downto 0);
    signal conv233_3794 : std_logic_vector(31 downto 0);
    signal conv24_3330 : std_logic_vector(31 downto 0);
    signal conv27_3343 : std_logic_vector(31 downto 0);
    signal conv2_3280 : std_logic_vector(15 downto 0);
    signal conv48_3361 : std_logic_vector(15 downto 0);
    signal conv4_3293 : std_logic_vector(15 downto 0);
    signal conv51_3374 : std_logic_vector(15 downto 0);
    signal conv60_3386 : std_logic_vector(15 downto 0);
    signal conv63_3399 : std_logic_vector(15 downto 0);
    signal conv82_3417 : std_logic_vector(15 downto 0);
    signal conv85_3430 : std_logic_vector(15 downto 0);
    signal conv91_3442 : std_logic_vector(15 downto 0);
    signal conv94_3455 : std_logic_vector(15 downto 0);
    signal conv98_3467 : std_logic_vector(31 downto 0);
    signal idxprom217_3743 : std_logic_vector(63 downto 0);
    signal idxprom_3720 : std_logic_vector(63 downto 0);
    signal inc241_3803 : std_logic_vector(15 downto 0);
    signal inc241x_xinput_dim0x_x2_3808 : std_logic_vector(15 downto 0);
    signal inc_3790 : std_logic_vector(15 downto 0);
    signal indvar_3620 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_3853 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_3841 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_3641 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_3835 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_3634 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_3815 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_3828 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_3627 : std_logic_vector(15 downto 0);
    signal mul185_3673 : std_logic_vector(15 downto 0);
    signal mul207_3695 : std_logic_vector(63 downto 0);
    signal mul209_3705 : std_logic_vector(63 downto 0);
    signal mul_3663 : std_logic_vector(15 downto 0);
    signal ptr_deref_3730_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3730_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3730_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3730_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3730_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3752_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3752_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3752_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3752_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3752_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3752_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl100_3473 : std_logic_vector(31 downto 0);
    signal shl105_3491 : std_logic_vector(31 downto 0);
    signal shl110_3509 : std_logic_vector(31 downto 0);
    signal shl132_3540 : std_logic_vector(63 downto 0);
    signal shl13_3311 : std_logic_vector(31 downto 0);
    signal shl144_3565 : std_logic_vector(63 downto 0);
    signal shl25_3336 : std_logic_vector(31 downto 0);
    signal shl49_3367 : std_logic_vector(15 downto 0);
    signal shl61_3392 : std_logic_vector(15 downto 0);
    signal shl83_3423 : std_logic_vector(15 downto 0);
    signal shl92_3448 : std_logic_vector(15 downto 0);
    signal shl_3286 : std_logic_vector(15 downto 0);
    signal shr157262_3590 : std_logic_vector(15 downto 0);
    signal shr212_3716 : std_logic_vector(31 downto 0);
    signal shr216_3737 : std_logic_vector(63 downto 0);
    signal shr261_3584 : std_logic_vector(15 downto 0);
    signal sub179_3668 : std_logic_vector(15 downto 0);
    signal sub192_3617 : std_logic_vector(15 downto 0);
    signal sub193_3678 : std_logic_vector(15 downto 0);
    signal sub_3606 : std_logic_vector(15 downto 0);
    signal tmp1_3653 : std_logic_vector(31 downto 0);
    signal tmp214_3731 : std_logic_vector(63 downto 0);
    signal type_cast_3284_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3309_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3334_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3365_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3390_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3421_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3446_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3471_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3489_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3507_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3538_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3563_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3582_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3588_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3599_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3610_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3624_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3626_wire : std_logic_vector(31 downto 0);
    signal type_cast_3631_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3633_wire : std_logic_vector(15 downto 0);
    signal type_cast_3638_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3640_wire : std_logic_vector(15 downto 0);
    signal type_cast_3644_wire : std_logic_vector(15 downto 0);
    signal type_cast_3646_wire : std_logic_vector(15 downto 0);
    signal type_cast_3651_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3714_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3735_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3741_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_3762_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3780_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3788_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3812_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3832_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3834_wire : std_logic_vector(15 downto 0);
    signal type_cast_3838_wire : std_logic_vector(15 downto 0);
    signal type_cast_3840_wire : std_logic_vector(15 downto 0);
    signal type_cast_3844_wire : std_logic_vector(15 downto 0);
    signal type_cast_3846_wire : std_logic_vector(15 downto 0);
    signal type_cast_3851_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3859_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_3725_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3725_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3725_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3725_resized_base_address <= "00000000000000";
    array_obj_ref_3748_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3748_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3748_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3748_resized_base_address <= "00000000000000";
    ptr_deref_3730_word_offset_0 <= "00000000000000";
    ptr_deref_3752_word_offset_0 <= "00000000000000";
    type_cast_3284_wire_constant <= "0000000000001000";
    type_cast_3309_wire_constant <= "00000000000000000000000000001000";
    type_cast_3334_wire_constant <= "00000000000000000000000000001000";
    type_cast_3365_wire_constant <= "0000000000001000";
    type_cast_3390_wire_constant <= "0000000000001000";
    type_cast_3421_wire_constant <= "0000000000001000";
    type_cast_3446_wire_constant <= "0000000000001000";
    type_cast_3471_wire_constant <= "00000000000000000000000000001000";
    type_cast_3489_wire_constant <= "00000000000000000000000000001000";
    type_cast_3507_wire_constant <= "00000000000000000000000000001000";
    type_cast_3538_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_3563_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_3582_wire_constant <= "0000000000000010";
    type_cast_3588_wire_constant <= "0000000000000001";
    type_cast_3599_wire_constant <= "1111111111111111";
    type_cast_3610_wire_constant <= "1111111111111111";
    type_cast_3624_wire_constant <= "00000000000000000000000000000000";
    type_cast_3631_wire_constant <= "0000000000000000";
    type_cast_3638_wire_constant <= "0000000000000000";
    type_cast_3651_wire_constant <= "00000000000000000000000000000100";
    type_cast_3714_wire_constant <= "00000000000000000000000000000010";
    type_cast_3735_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_3741_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_3762_wire_constant <= "00000000000000000000000000000100";
    type_cast_3780_wire_constant <= "0000000000000100";
    type_cast_3788_wire_constant <= "0000000000000001";
    type_cast_3812_wire_constant <= "0000000000000000";
    type_cast_3832_wire_constant <= "0000000000000000";
    type_cast_3851_wire_constant <= "00000000000000000000000000000001";
    type_cast_3859_wire_constant <= "00000001";
    phi_stmt_3620: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3624_wire_constant & type_cast_3626_wire;
      req <= phi_stmt_3620_req_0 & phi_stmt_3620_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3620",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3620_ack_0,
          idata => idata,
          odata => indvar_3620,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3620
    phi_stmt_3627: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3631_wire_constant & type_cast_3633_wire;
      req <= phi_stmt_3627_req_0 & phi_stmt_3627_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3627",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3627_ack_0,
          idata => idata,
          odata => input_dim2x_x1_3627,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3627
    phi_stmt_3634: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3638_wire_constant & type_cast_3640_wire;
      req <= phi_stmt_3634_req_0 & phi_stmt_3634_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3634",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3634_ack_0,
          idata => idata,
          odata => input_dim1x_x1_3634,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3634
    phi_stmt_3641: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3644_wire & type_cast_3646_wire;
      req <= phi_stmt_3641_req_0 & phi_stmt_3641_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3641",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3641_ack_0,
          idata => idata,
          odata => input_dim0x_x2_3641,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3641
    phi_stmt_3828: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3832_wire_constant & type_cast_3834_wire;
      req <= phi_stmt_3828_req_0 & phi_stmt_3828_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3828",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3828_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_3828,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3828
    phi_stmt_3835: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3838_wire & type_cast_3840_wire;
      req <= phi_stmt_3835_req_0 & phi_stmt_3835_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3835",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3835_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_3835,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3835
    phi_stmt_3841: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3844_wire & type_cast_3846_wire;
      req <= phi_stmt_3841_req_0 & phi_stmt_3841_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3841",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3841_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_3841,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3841
    -- flow-through select operator MUX_3814_inst
    input_dim1x_x2_3815 <= type_cast_3812_wire_constant when (cmp237_3799(0) /=  '0') else inc_3790;
    addr_of_3726_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3726_final_reg_req_0;
      addr_of_3726_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3726_final_reg_req_1;
      addr_of_3726_final_reg_ack_1<= rack(0);
      addr_of_3726_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3726_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3725_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx213_3727,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3749_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3749_final_reg_req_0;
      addr_of_3749_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3749_final_reg_req_1;
      addr_of_3749_final_reg_ack_1<= rack(0);
      addr_of_3749_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3749_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3748_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx218_3750,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3279_inst_req_0;
      type_cast_3279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3279_inst_req_1;
      type_cast_3279_inst_ack_1<= rack(0);
      type_cast_3279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_3276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_3280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3292_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3292_inst_req_0;
      type_cast_3292_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3292_inst_req_1;
      type_cast_3292_inst_ack_1<= rack(0);
      type_cast_3292_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3292_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_3289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_3293,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3304_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3304_inst_req_0;
      type_cast_3304_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3304_inst_req_1;
      type_cast_3304_inst_ack_1<= rack(0);
      type_cast_3304_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3304_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call7_3301,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_3305,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3317_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3317_inst_req_0;
      type_cast_3317_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3317_inst_req_1;
      type_cast_3317_inst_ack_1<= rack(0);
      type_cast_3317_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3317_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_3314,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_3318,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3329_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3329_inst_req_0;
      type_cast_3329_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3329_inst_req_1;
      type_cast_3329_inst_ack_1<= rack(0);
      type_cast_3329_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3329_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_3326,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_3330,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3342_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3342_inst_req_0;
      type_cast_3342_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3342_inst_req_1;
      type_cast_3342_inst_ack_1<= rack(0);
      type_cast_3342_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3342_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_3339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_3343,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3360_inst_req_0;
      type_cast_3360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3360_inst_req_1;
      type_cast_3360_inst_ack_1<= rack(0);
      type_cast_3360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call43_3357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_3361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3373_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3373_inst_req_0;
      type_cast_3373_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3373_inst_req_1;
      type_cast_3373_inst_ack_1<= rack(0);
      type_cast_3373_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3373_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_3370,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_3374,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3385_inst_req_0;
      type_cast_3385_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3385_inst_req_1;
      type_cast_3385_inst_ack_1<= rack(0);
      type_cast_3385_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3385_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_3382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_3386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3398_inst_req_0;
      type_cast_3398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3398_inst_req_1;
      type_cast_3398_inst_ack_1<= rack(0);
      type_cast_3398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call62_3395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_3399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3416_inst_req_0;
      type_cast_3416_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3416_inst_req_1;
      type_cast_3416_inst_ack_1<= rack(0);
      type_cast_3416_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3416_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call79_3413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_3417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3429_inst_req_0;
      type_cast_3429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3429_inst_req_1;
      type_cast_3429_inst_ack_1<= rack(0);
      type_cast_3429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call84_3426,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_3430,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3441_inst_req_0;
      type_cast_3441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3441_inst_req_1;
      type_cast_3441_inst_ack_1<= rack(0);
      type_cast_3441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_3438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_3442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3454_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3454_inst_req_0;
      type_cast_3454_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3454_inst_req_1;
      type_cast_3454_inst_ack_1<= rack(0);
      type_cast_3454_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3454_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_3451,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_3455,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3466_inst_req_0;
      type_cast_3466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3466_inst_req_1;
      type_cast_3466_inst_ack_1<= rack(0);
      type_cast_3466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_3463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_3467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3479_inst_req_0;
      type_cast_3479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3479_inst_req_1;
      type_cast_3479_inst_ack_1<= rack(0);
      type_cast_3479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_3476,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv102_3480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3497_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3497_inst_req_0;
      type_cast_3497_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3497_inst_req_1;
      type_cast_3497_inst_ack_1<= rack(0);
      type_cast_3497_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3497_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_3494,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_3498,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3515_inst_req_0;
      type_cast_3515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3515_inst_req_1;
      type_cast_3515_inst_ack_1<= rack(0);
      type_cast_3515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_3512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_3516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3533_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3533_inst_req_0;
      type_cast_3533_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3533_inst_req_1;
      type_cast_3533_inst_ack_1<= rack(0);
      type_cast_3533_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3533_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call126_3530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_3534,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3546_inst_req_0;
      type_cast_3546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3546_inst_req_1;
      type_cast_3546_inst_ack_1<= rack(0);
      type_cast_3546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3546_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_3543,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_3547,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3558_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3558_inst_req_0;
      type_cast_3558_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3558_inst_req_1;
      type_cast_3558_inst_ack_1<= rack(0);
      type_cast_3558_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3558_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call138_3555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_3559,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3571_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3571_inst_req_0;
      type_cast_3571_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3571_inst_req_1;
      type_cast_3571_inst_ack_1<= rack(0);
      type_cast_3571_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3571_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_3568,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv146_3572,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3626_inst_req_0;
      type_cast_3626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3626_inst_req_1;
      type_cast_3626_inst_ack_1<= rack(0);
      type_cast_3626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_3853,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3626_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3633_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3633_inst_req_0;
      type_cast_3633_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3633_inst_req_1;
      type_cast_3633_inst_ack_1<= rack(0);
      type_cast_3633_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3633_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_3828,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3633_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3640_inst_req_0;
      type_cast_3640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3640_inst_req_1;
      type_cast_3640_inst_ack_1<= rack(0);
      type_cast_3640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_3835,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3640_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3644_inst_req_0;
      type_cast_3644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3644_inst_req_1;
      type_cast_3644_inst_ack_1<= rack(0);
      type_cast_3644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_3841,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3644_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3646_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3646_inst_req_0;
      type_cast_3646_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3646_inst_req_1;
      type_cast_3646_inst_ack_1<= rack(0);
      type_cast_3646_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3646_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add158_3595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3646_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3681_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3681_inst_req_0;
      type_cast_3681_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3681_inst_req_1;
      type_cast_3681_inst_ack_1<= rack(0);
      type_cast_3681_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3681_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_3627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv196_3682,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3685_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3685_inst_req_0;
      type_cast_3685_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3685_inst_req_1;
      type_cast_3685_inst_ack_1<= rack(0);
      type_cast_3685_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3685_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub193_3678,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv201_3686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3689_inst_req_0;
      type_cast_3689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3689_inst_req_1;
      type_cast_3689_inst_ack_1<= rack(0);
      type_cast_3689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub179_3668,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_3690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3719_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3719_inst_req_0;
      type_cast_3719_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3719_inst_req_1;
      type_cast_3719_inst_ack_1<= rack(0);
      type_cast_3719_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3719_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr212_3716,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3720,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3757_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3757_inst_req_0;
      type_cast_3757_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3757_inst_req_1;
      type_cast_3757_inst_ack_1<= rack(0);
      type_cast_3757_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3757_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_3627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv221_3758,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3793_inst_req_0;
      type_cast_3793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3793_inst_req_1;
      type_cast_3793_inst_ack_1<= rack(0);
      type_cast_3793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_3790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv233_3794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3802_inst_req_0;
      type_cast_3802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3802_inst_req_1;
      type_cast_3802_inst_ack_1<= rack(0);
      type_cast_3802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp237_3799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc241_3803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3834_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3834_inst_req_0;
      type_cast_3834_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3834_inst_req_1;
      type_cast_3834_inst_ack_1<= rack(0);
      type_cast_3834_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3834_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add229_3782,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3834_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3838_inst_req_0;
      type_cast_3838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3838_inst_req_1;
      type_cast_3838_inst_ack_1<= rack(0);
      type_cast_3838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_3634,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3838_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3840_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3840_inst_req_0;
      type_cast_3840_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3840_inst_req_1;
      type_cast_3840_inst_ack_1<= rack(0);
      type_cast_3840_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3840_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_3815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3840_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3844_inst_req_0;
      type_cast_3844_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3844_inst_req_1;
      type_cast_3844_inst_ack_1<= rack(0);
      type_cast_3844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_3641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3844_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3846_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3846_inst_req_0;
      type_cast_3846_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3846_inst_req_1;
      type_cast_3846_inst_ack_1<= rack(0);
      type_cast_3846_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3846_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc241x_xinput_dim0x_x2_3808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3846_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_3725_index_1_rename
    process(R_idxprom_3724_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3724_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3724_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3725_index_1_resize
    process(idxprom_3720) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3720;
      ov := iv(13 downto 0);
      R_idxprom_3724_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3725_root_address_inst
    process(array_obj_ref_3725_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3725_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3725_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3748_index_1_rename
    process(R_idxprom217_3747_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom217_3747_resized;
      ov(13 downto 0) := iv;
      R_idxprom217_3747_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3748_index_1_resize
    process(idxprom217_3743) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom217_3743;
      ov := iv(13 downto 0);
      R_idxprom217_3747_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3748_root_address_inst
    process(array_obj_ref_3748_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3748_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3748_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3730_addr_0
    process(ptr_deref_3730_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3730_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3730_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3730_base_resize
    process(arrayidx213_3727) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx213_3727;
      ov := iv(13 downto 0);
      ptr_deref_3730_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3730_gather_scatter
    process(ptr_deref_3730_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3730_data_0;
      ov(63 downto 0) := iv;
      tmp214_3731 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3730_root_address_inst
    process(ptr_deref_3730_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3730_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3730_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3752_addr_0
    process(ptr_deref_3752_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3752_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3752_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3752_base_resize
    process(arrayidx218_3750) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx218_3750;
      ov := iv(13 downto 0);
      ptr_deref_3752_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3752_gather_scatter
    process(tmp214_3731) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp214_3731;
      ov(63 downto 0) := iv;
      ptr_deref_3752_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3752_root_address_inst
    process(ptr_deref_3752_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3752_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3752_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3770_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_3769;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3770_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3770_branch_req_0,
          ack0 => if_stmt_3770_branch_ack_0,
          ack1 => if_stmt_3770_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3821_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp247_3820;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3821_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3821_branch_req_0,
          ack0 => if_stmt_3821_branch_ack_0,
          ack1 => if_stmt_3821_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3594_inst
    process(shr261_3584, shr157262_3590) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr261_3584, shr157262_3590, tmp_var);
      add158_3595 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3600_inst
    process(add52_3379) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add52_3379, type_cast_3599_wire_constant, tmp_var);
      add176_3601 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3611_inst
    process(add64_3404) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add64_3404, type_cast_3610_wire_constant, tmp_var);
      add189_3612 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3667_inst
    process(sub_3606, mul_3663) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_3606, mul_3663, tmp_var);
      sub179_3668 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3677_inst
    process(sub192_3617, mul185_3673) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub192_3617, mul185_3673, tmp_var);
      sub193_3678 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3781_inst
    process(input_dim2x_x1_3627) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_3627, type_cast_3780_wire_constant, tmp_var);
      add229_3782 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3789_inst
    process(input_dim1x_x1_3634) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_3634, type_cast_3788_wire_constant, tmp_var);
      inc_3790 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3807_inst
    process(inc241_3803, input_dim0x_x2_3641) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc241_3803, input_dim0x_x2_3641, tmp_var);
      inc241x_xinput_dim0x_x2_3808 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3657_inst
    process(add113_3521, tmp1_3653) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add113_3521, tmp1_3653, tmp_var);
      add_src_0x_x0_3658 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3763_inst
    process(conv221_3758) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv221_3758, type_cast_3762_wire_constant, tmp_var);
      add222_3764 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3852_inst
    process(indvar_3620) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_3620, type_cast_3851_wire_constant, tmp_var);
      indvarx_xnext_3853 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_3699_inst
    process(mul207_3695, conv201_3686) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul207_3695, conv201_3686, tmp_var);
      add208_3700 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_3709_inst
    process(mul209_3705, conv196_3682) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul209_3705, conv196_3682, tmp_var);
      add210_3710 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_3742_inst
    process(shr216_3737) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr216_3737, type_cast_3741_wire_constant, tmp_var);
      idxprom217_3743 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_3819_inst
    process(inc241x_xinput_dim0x_x2_3808, add_3298) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc241x_xinput_dim0x_x2_3808, add_3298, tmp_var);
      cmp247_3820 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3798_inst
    process(conv233_3794, add16_3323) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv233_3794, add16_3323, tmp_var);
      cmp237_3799 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3583_inst
    process(add_3298) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_3298, type_cast_3582_wire_constant, tmp_var);
      shr261_3584 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_3589_inst
    process(add_3298) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_3298, type_cast_3588_wire_constant, tmp_var);
      shr157262_3590 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3715_inst
    process(add_src_0x_x0_3658) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_3658, type_cast_3714_wire_constant, tmp_var);
      shr212_3716 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_3736_inst
    process(add210_3710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add210_3710, type_cast_3735_wire_constant, tmp_var);
      shr216_3737 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3662_inst
    process(input_dim0x_x2_3641, add86_3435) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_3641, add86_3435, tmp_var);
      mul_3663 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3672_inst
    process(input_dim1x_x1_3634, add86_3435) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_3634, add86_3435, tmp_var);
      mul185_3673 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3652_inst
    process(indvar_3620) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_3620, type_cast_3651_wire_constant, tmp_var);
      tmp1_3653 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_3694_inst
    process(conv206_3690, add135_3552) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv206_3690, add135_3552, tmp_var);
      mul207_3695 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_3704_inst
    process(add208_3700, add147_3577) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add208_3700, add147_3577, tmp_var);
      mul209_3705 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_3297_inst
    process(shl_3286, conv4_3293) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_3286, conv4_3293, tmp_var);
      add_3298 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_3378_inst
    process(shl49_3367, conv51_3374) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl49_3367, conv51_3374, tmp_var);
      add52_3379 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_3403_inst
    process(shl61_3392, conv63_3399) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl61_3392, conv63_3399, tmp_var);
      add64_3404 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_3434_inst
    process(shl83_3423, conv85_3430) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl83_3423, conv85_3430, tmp_var);
      add86_3435 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_3459_inst
    process(shl92_3448, conv94_3455) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_3448, conv94_3455, tmp_var);
      add95_3460 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_3322_inst
    process(shl13_3311, conv15_3318) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl13_3311, conv15_3318, tmp_var);
      add16_3323 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_3347_inst
    process(shl25_3336, conv27_3343) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl25_3336, conv27_3343, tmp_var);
      add28_3348 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_3484_inst
    process(shl100_3473, conv102_3480) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_3473, conv102_3480, tmp_var);
      add103_3485 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_3502_inst
    process(shl105_3491, conv107_3498) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_3491, conv107_3498, tmp_var);
      add108_3503 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_3520_inst
    process(shl110_3509, conv112_3516) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_3509, conv112_3516, tmp_var);
      add113_3521 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_3551_inst
    process(shl132_3540, conv134_3547) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_3540, conv134_3547, tmp_var);
      add135_3552 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_3576_inst
    process(shl144_3565, conv146_3572) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_3565, conv146_3572, tmp_var);
      add147_3577 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_3285_inst
    process(conv2_3280) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv2_3280, type_cast_3284_wire_constant, tmp_var);
      shl_3286 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_3366_inst
    process(conv48_3361) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv48_3361, type_cast_3365_wire_constant, tmp_var);
      shl49_3367 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_3391_inst
    process(conv60_3386) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv60_3386, type_cast_3390_wire_constant, tmp_var);
      shl61_3392 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_3422_inst
    process(conv82_3417) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv82_3417, type_cast_3421_wire_constant, tmp_var);
      shl83_3423 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_3447_inst
    process(conv91_3442) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_3442, type_cast_3446_wire_constant, tmp_var);
      shl92_3448 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3310_inst
    process(conv12_3305) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv12_3305, type_cast_3309_wire_constant, tmp_var);
      shl13_3311 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3335_inst
    process(conv24_3330) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv24_3330, type_cast_3334_wire_constant, tmp_var);
      shl25_3336 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3472_inst
    process(conv98_3467) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv98_3467, type_cast_3471_wire_constant, tmp_var);
      shl100_3473 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3490_inst
    process(add103_3485) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add103_3485, type_cast_3489_wire_constant, tmp_var);
      shl105_3491 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3508_inst
    process(add108_3503) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_3503, type_cast_3507_wire_constant, tmp_var);
      shl110_3509 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_3539_inst
    process(conv131_3534) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_3534, type_cast_3538_wire_constant, tmp_var);
      shl132_3540 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_3564_inst
    process(conv143_3559) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv143_3559, type_cast_3563_wire_constant, tmp_var);
      shl144_3565 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_3605_inst
    process(add176_3601, add95_3460) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add176_3601, add95_3460, tmp_var);
      sub_3606 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_3616_inst
    process(add189_3612, add95_3460) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add189_3612, add95_3460, tmp_var);
      sub192_3617 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_3768_inst
    process(add222_3764, add28_3348) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add222_3764, add28_3348, tmp_var);
      cmp_3769 <= tmp_var; --
    end process;
    -- shared split operator group (52) : array_obj_ref_3725_index_offset 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3724_scaled;
      array_obj_ref_3725_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3725_index_offset_req_0;
      array_obj_ref_3725_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3725_index_offset_req_1;
      array_obj_ref_3725_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : array_obj_ref_3748_index_offset 
    ApIntAdd_group_53: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom217_3747_scaled;
      array_obj_ref_3748_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3748_index_offset_req_0;
      array_obj_ref_3748_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3748_index_offset_req_1;
      array_obj_ref_3748_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_53_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_53_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_53",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared load operator group (0) : ptr_deref_3730_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3730_load_0_req_0;
      ptr_deref_3730_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3730_load_0_req_1;
      ptr_deref_3730_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3730_word_address_0;
      ptr_deref_3730_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3752_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3752_store_0_req_0;
      ptr_deref_3752_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3752_store_0_req_1;
      ptr_deref_3752_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3752_word_address_0;
      data_in <= ptr_deref_3752_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_3450_inst RPIPE_Block3_start_3350_inst RPIPE_Block3_start_3353_inst RPIPE_Block3_start_3462_inst RPIPE_Block3_start_3356_inst RPIPE_Block3_start_3369_inst RPIPE_Block3_start_3425_inst RPIPE_Block3_start_3437_inst RPIPE_Block3_start_3338_inst RPIPE_Block3_start_3567_inst RPIPE_Block3_start_3554_inst RPIPE_Block3_start_3542_inst RPIPE_Block3_start_3412_inst RPIPE_Block3_start_3325_inst RPIPE_Block3_start_3409_inst RPIPE_Block3_start_3313_inst RPIPE_Block3_start_3529_inst RPIPE_Block3_start_3406_inst RPIPE_Block3_start_3526_inst RPIPE_Block3_start_3523_inst RPIPE_Block3_start_3511_inst RPIPE_Block3_start_3394_inst RPIPE_Block3_start_3300_inst RPIPE_Block3_start_3381_inst RPIPE_Block3_start_3493_inst RPIPE_Block3_start_3288_inst RPIPE_Block3_start_3475_inst RPIPE_Block3_start_3275_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 27 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 27 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant outBUFs : IntegerArray(27 downto 0) := (27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      reqL_unguarded(27) <= RPIPE_Block3_start_3450_inst_req_0;
      reqL_unguarded(26) <= RPIPE_Block3_start_3350_inst_req_0;
      reqL_unguarded(25) <= RPIPE_Block3_start_3353_inst_req_0;
      reqL_unguarded(24) <= RPIPE_Block3_start_3462_inst_req_0;
      reqL_unguarded(23) <= RPIPE_Block3_start_3356_inst_req_0;
      reqL_unguarded(22) <= RPIPE_Block3_start_3369_inst_req_0;
      reqL_unguarded(21) <= RPIPE_Block3_start_3425_inst_req_0;
      reqL_unguarded(20) <= RPIPE_Block3_start_3437_inst_req_0;
      reqL_unguarded(19) <= RPIPE_Block3_start_3338_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Block3_start_3567_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Block3_start_3554_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Block3_start_3542_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Block3_start_3412_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Block3_start_3325_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Block3_start_3409_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_3313_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_3529_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_3406_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_3526_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_3523_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_3511_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_3394_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_3300_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_3381_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_3493_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_3288_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_3475_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_3275_inst_req_0;
      RPIPE_Block3_start_3450_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_Block3_start_3350_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_Block3_start_3353_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_Block3_start_3462_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_Block3_start_3356_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_Block3_start_3369_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_Block3_start_3425_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_Block3_start_3437_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_Block3_start_3338_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Block3_start_3567_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Block3_start_3554_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Block3_start_3542_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Block3_start_3412_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Block3_start_3325_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Block3_start_3409_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_3313_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_3529_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_3406_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_3526_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_3523_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_3511_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_3394_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_3300_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_3381_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_3493_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_3288_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_3475_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_3275_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(27) <= RPIPE_Block3_start_3450_inst_req_1;
      reqR_unguarded(26) <= RPIPE_Block3_start_3350_inst_req_1;
      reqR_unguarded(25) <= RPIPE_Block3_start_3353_inst_req_1;
      reqR_unguarded(24) <= RPIPE_Block3_start_3462_inst_req_1;
      reqR_unguarded(23) <= RPIPE_Block3_start_3356_inst_req_1;
      reqR_unguarded(22) <= RPIPE_Block3_start_3369_inst_req_1;
      reqR_unguarded(21) <= RPIPE_Block3_start_3425_inst_req_1;
      reqR_unguarded(20) <= RPIPE_Block3_start_3437_inst_req_1;
      reqR_unguarded(19) <= RPIPE_Block3_start_3338_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Block3_start_3567_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Block3_start_3554_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Block3_start_3542_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Block3_start_3412_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Block3_start_3325_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Block3_start_3409_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_3313_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_3529_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_3406_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_3526_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_3523_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_3511_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_3394_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_3300_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_3381_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_3493_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_3288_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_3475_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_3275_inst_req_1;
      RPIPE_Block3_start_3450_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_Block3_start_3350_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_Block3_start_3353_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_Block3_start_3462_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_Block3_start_3356_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_Block3_start_3369_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_Block3_start_3425_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_Block3_start_3437_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_Block3_start_3338_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Block3_start_3567_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Block3_start_3554_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Block3_start_3542_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Block3_start_3412_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Block3_start_3325_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Block3_start_3409_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_3313_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_3529_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_3406_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_3526_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_3523_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_3511_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_3394_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_3300_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_3381_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_3493_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_3288_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_3475_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_3275_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      call93_3451 <= data_out(223 downto 216);
      call31_3351 <= data_out(215 downto 208);
      call38_3354 <= data_out(207 downto 200);
      call97_3463 <= data_out(199 downto 192);
      call43_3357 <= data_out(191 downto 184);
      call50_3370 <= data_out(183 downto 176);
      call84_3426 <= data_out(175 downto 168);
      call88_3438 <= data_out(167 downto 160);
      call26_3339 <= data_out(159 downto 152);
      call145_3568 <= data_out(151 downto 144);
      call138_3555 <= data_out(143 downto 136);
      call133_3543 <= data_out(135 downto 128);
      call79_3413 <= data_out(127 downto 120);
      call19_3326 <= data_out(119 downto 112);
      call74_3410 <= data_out(111 downto 104);
      call14_3314 <= data_out(103 downto 96);
      call126_3530 <= data_out(95 downto 88);
      call67_3407 <= data_out(87 downto 80);
      call121_3527 <= data_out(79 downto 72);
      call114_3524 <= data_out(71 downto 64);
      call111_3512 <= data_out(63 downto 56);
      call62_3395 <= data_out(55 downto 48);
      call7_3301 <= data_out(47 downto 40);
      call55_3382 <= data_out(39 downto 32);
      call106_3494 <= data_out(31 downto 24);
      call3_3289 <= data_out(23 downto 16);
      call101_3476 <= data_out(15 downto 8);
      call_3276 <= data_out(7 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 8,  num_reqs => 28,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_3857_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_3857_inst_req_0;
      WPIPE_Block3_done_3857_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_3857_inst_req_1;
      WPIPE_Block3_done_3857_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_3859_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_28_load_0_req_0 : boolean;
  signal LOAD_count_28_load_0_ack_0 : boolean;
  signal LOAD_count_28_load_0_req_1 : boolean;
  signal LOAD_count_28_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_29/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_sample_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_update_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$entry
      -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_1); -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_sample_completed_
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$exit
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_req
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_29/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_update_completed_
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_ack
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_28_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_28_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_28_word_address_0 <= "0";
    -- equivalence LOAD_count_28_gather_scatter
    process(LOAD_count_28_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_28_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_28_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_28_load_0_req_0;
      LOAD_count_28_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_28_load_0_req_1;
      LOAD_count_28_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_28_word_address_0;
      LOAD_count_28_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(7 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(7 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(7 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(7 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(7 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(7 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(7 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(7 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(7 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(7 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(7 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(7 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(7 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(7 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(7 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(7 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(7 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
