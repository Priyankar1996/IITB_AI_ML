-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    row_in : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
    input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe4_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 48)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal row_in_buffer :  std_logic_vector(15 downto 0);
  signal row_in_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal W_fetch_val2_322_delayed_13_0_340_inst_req_1 : boolean;
  signal W_fetch_val2_322_delayed_13_0_340_inst_ack_0 : boolean;
  signal W_fetch_val2_322_delayed_13_0_340_inst_req_0 : boolean;
  signal W_fn2_320_delayed_13_0_337_inst_req_1 : boolean;
  signal type_cast_371_inst_req_0 : boolean;
  signal W_fetch_val2_322_delayed_13_0_340_inst_ack_1 : boolean;
  signal addr_of_327_final_reg_ack_1 : boolean;
  signal array_obj_ref_326_index_offset_ack_0 : boolean;
  signal ptr_deref_335_load_0_ack_1 : boolean;
  signal array_obj_ref_326_index_offset_req_0 : boolean;
  signal ptr_deref_263_load_0_ack_1 : boolean;
  signal ptr_deref_52_load_0_req_0 : boolean;
  signal ptr_deref_52_load_0_ack_0 : boolean;
  signal ptr_deref_263_load_0_req_1 : boolean;
  signal ptr_deref_52_load_0_req_1 : boolean;
  signal ptr_deref_52_load_0_ack_1 : boolean;
  signal type_cast_299_inst_ack_1 : boolean;
  signal array_obj_ref_75_index_offset_req_0 : boolean;
  signal array_obj_ref_75_index_offset_ack_0 : boolean;
  signal addr_of_327_final_reg_req_1 : boolean;
  signal ptr_deref_335_load_0_req_1 : boolean;
  signal array_obj_ref_61_index_offset_req_0 : boolean;
  signal array_obj_ref_61_index_offset_ack_0 : boolean;
  signal W_fn2_320_delayed_13_0_337_inst_ack_0 : boolean;
  signal array_obj_ref_61_index_offset_req_1 : boolean;
  signal array_obj_ref_61_index_offset_ack_1 : boolean;
  signal W_fn2_314_delayed_7_0_329_inst_ack_0 : boolean;
  signal W_fn2_320_delayed_13_0_337_inst_req_0 : boolean;
  signal addr_of_62_final_reg_req_0 : boolean;
  signal addr_of_62_final_reg_ack_0 : boolean;
  signal addr_of_62_final_reg_req_1 : boolean;
  signal addr_of_62_final_reg_ack_1 : boolean;
  signal ptr_deref_335_load_0_ack_0 : boolean;
  signal addr_of_327_final_reg_ack_0 : boolean;
  signal addr_of_327_final_reg_req_0 : boolean;
  signal ptr_deref_66_load_0_req_0 : boolean;
  signal ptr_deref_66_load_0_ack_0 : boolean;
  signal ptr_deref_66_load_0_req_1 : boolean;
  signal ptr_deref_66_load_0_ack_1 : boolean;
  signal ptr_deref_335_load_0_req_0 : boolean;
  signal phi_stmt_102_ack_0 : boolean;
  signal array_obj_ref_75_index_offset_req_1 : boolean;
  signal array_obj_ref_75_index_offset_ack_1 : boolean;
  signal W_fn2_314_delayed_7_0_329_inst_req_0 : boolean;
  signal addr_of_76_final_reg_req_0 : boolean;
  signal addr_of_76_final_reg_ack_0 : boolean;
  signal addr_of_76_final_reg_req_1 : boolean;
  signal addr_of_76_final_reg_ack_1 : boolean;
  signal addr_of_255_final_reg_ack_0 : boolean;
  signal type_cast_299_inst_req_1 : boolean;
  signal ptr_deref_263_load_0_ack_0 : boolean;
  signal ptr_deref_80_load_0_req_0 : boolean;
  signal ptr_deref_80_load_0_ack_0 : boolean;
  signal addr_of_255_final_reg_ack_1 : boolean;
  signal ptr_deref_263_load_0_req_0 : boolean;
  signal ptr_deref_80_load_0_req_1 : boolean;
  signal ptr_deref_80_load_0_ack_1 : boolean;
  signal type_cast_299_inst_ack_0 : boolean;
  signal type_cast_299_inst_req_0 : boolean;
  signal array_obj_ref_93_index_offset_req_0 : boolean;
  signal array_obj_ref_93_index_offset_ack_0 : boolean;
  signal array_obj_ref_93_index_offset_req_1 : boolean;
  signal array_obj_ref_93_index_offset_ack_1 : boolean;
  signal addr_of_94_final_reg_req_0 : boolean;
  signal addr_of_94_final_reg_ack_0 : boolean;
  signal addr_of_94_final_reg_req_1 : boolean;
  signal addr_of_94_final_reg_ack_1 : boolean;
  signal ptr_deref_98_load_0_req_0 : boolean;
  signal ptr_deref_98_load_0_ack_0 : boolean;
  signal addr_of_255_final_reg_req_1 : boolean;
  signal ptr_deref_98_load_0_req_1 : boolean;
  signal ptr_deref_98_load_0_ack_1 : boolean;
  signal W_fn2_320_delayed_13_0_337_inst_ack_1 : boolean;
  signal array_obj_ref_326_index_offset_ack_1 : boolean;
  signal do_while_stmt_100_branch_req_0 : boolean;
  signal array_obj_ref_326_index_offset_req_1 : boolean;
  signal addr_of_255_final_reg_req_0 : boolean;
  signal phi_stmt_102_req_1 : boolean;
  signal phi_stmt_102_req_0 : boolean;
  signal n_fetch_val1_276_132_buf_req_0 : boolean;
  signal n_fetch_val1_276_132_buf_ack_0 : boolean;
  signal n_fetch_val1_276_132_buf_req_1 : boolean;
  signal n_fetch_val1_276_132_buf_ack_1 : boolean;
  signal n_address1_236_106_buf_req_0 : boolean;
  signal n_address1_236_106_buf_ack_0 : boolean;
  signal n_address1_236_106_buf_req_1 : boolean;
  signal n_address1_236_106_buf_ack_1 : boolean;
  signal phi_stmt_107_req_1 : boolean;
  signal phi_stmt_107_req_0 : boolean;
  signal phi_stmt_107_ack_0 : boolean;
  signal type_cast_110_inst_req_0 : boolean;
  signal type_cast_110_inst_ack_0 : boolean;
  signal type_cast_110_inst_req_1 : boolean;
  signal type_cast_110_inst_ack_1 : boolean;
  signal W_fetch_val1_262_delayed_13_0_268_inst_ack_1 : boolean;
  signal W_fetch_val1_262_delayed_13_0_268_inst_req_1 : boolean;
  signal n_address2_308_111_buf_req_0 : boolean;
  signal n_address2_308_111_buf_ack_0 : boolean;
  signal n_address2_308_111_buf_req_1 : boolean;
  signal n_address2_308_111_buf_ack_1 : boolean;
  signal W_fetch_val1_262_delayed_13_0_268_inst_ack_0 : boolean;
  signal W_fetch_val1_262_delayed_13_0_268_inst_req_0 : boolean;
  signal phi_stmt_112_req_1 : boolean;
  signal phi_stmt_112_req_0 : boolean;
  signal phi_stmt_112_ack_0 : boolean;
  signal type_cast_115_inst_req_0 : boolean;
  signal type_cast_115_inst_ack_0 : boolean;
  signal type_cast_115_inst_req_1 : boolean;
  signal type_cast_115_inst_ack_1 : boolean;
  signal n_address3_380_116_buf_req_0 : boolean;
  signal n_address3_380_116_buf_ack_0 : boolean;
  signal W_fn1_254_delayed_7_0_257_inst_ack_1 : boolean;
  signal W_fn1_254_delayed_7_0_257_inst_req_1 : boolean;
  signal n_address3_380_116_buf_req_1 : boolean;
  signal n_address3_380_116_buf_ack_1 : boolean;
  signal phi_stmt_117_req_1 : boolean;
  signal phi_stmt_117_req_0 : boolean;
  signal phi_stmt_117_ack_0 : boolean;
  signal W_fn1_260_delayed_13_0_265_inst_ack_1 : boolean;
  signal W_fn1_260_delayed_13_0_265_inst_req_1 : boolean;
  signal type_cast_122_inst_req_0 : boolean;
  signal type_cast_122_inst_ack_0 : boolean;
  signal W_fn2_314_delayed_7_0_329_inst_ack_1 : boolean;
  signal type_cast_122_inst_req_1 : boolean;
  signal type_cast_122_inst_ack_1 : boolean;
  signal W_fn1_254_delayed_7_0_257_inst_ack_0 : boolean;
  signal W_fn1_254_delayed_7_0_257_inst_req_0 : boolean;
  signal W_fn1_260_delayed_13_0_265_inst_ack_0 : boolean;
  signal W_fn1_260_delayed_13_0_265_inst_req_0 : boolean;
  signal W_fn2_314_delayed_7_0_329_inst_req_1 : boolean;
  signal n_address4_452_123_buf_req_0 : boolean;
  signal n_address4_452_123_buf_ack_0 : boolean;
  signal n_address4_452_123_buf_req_1 : boolean;
  signal n_address4_452_123_buf_ack_1 : boolean;
  signal phi_stmt_124_req_1 : boolean;
  signal phi_stmt_124_req_0 : boolean;
  signal phi_stmt_124_ack_0 : boolean;
  signal n_mycounter_168_128_buf_req_0 : boolean;
  signal n_mycounter_168_128_buf_ack_0 : boolean;
  signal n_mycounter_168_128_buf_req_1 : boolean;
  signal n_mycounter_168_128_buf_ack_1 : boolean;
  signal phi_stmt_129_req_1 : boolean;
  signal phi_stmt_129_req_0 : boolean;
  signal phi_stmt_129_ack_0 : boolean;
  signal my_fetch1_53_131_buf_req_0 : boolean;
  signal my_fetch1_53_131_buf_ack_0 : boolean;
  signal my_fetch1_53_131_buf_req_1 : boolean;
  signal my_fetch1_53_131_buf_ack_1 : boolean;
  signal phi_stmt_133_req_1 : boolean;
  signal phi_stmt_133_req_0 : boolean;
  signal phi_stmt_133_ack_0 : boolean;
  signal my_fetch2_67_135_buf_req_0 : boolean;
  signal my_fetch2_67_135_buf_ack_0 : boolean;
  signal my_fetch2_67_135_buf_req_1 : boolean;
  signal my_fetch2_67_135_buf_ack_1 : boolean;
  signal type_cast_371_inst_ack_0 : boolean;
  signal type_cast_371_inst_req_1 : boolean;
  signal n_fetch_val2_348_136_buf_req_0 : boolean;
  signal n_fetch_val2_348_136_buf_ack_0 : boolean;
  signal n_fetch_val2_348_136_buf_req_1 : boolean;
  signal n_fetch_val2_348_136_buf_ack_1 : boolean;
  signal phi_stmt_137_req_1 : boolean;
  signal phi_stmt_137_req_0 : boolean;
  signal phi_stmt_137_ack_0 : boolean;
  signal my_fetch3_81_139_buf_req_0 : boolean;
  signal my_fetch3_81_139_buf_ack_0 : boolean;
  signal my_fetch3_81_139_buf_req_1 : boolean;
  signal my_fetch3_81_139_buf_ack_1 : boolean;
  signal n_fetch_val3_420_140_buf_req_0 : boolean;
  signal n_fetch_val3_420_140_buf_ack_0 : boolean;
  signal n_fetch_val3_420_140_buf_req_1 : boolean;
  signal n_fetch_val3_420_140_buf_ack_1 : boolean;
  signal phi_stmt_141_req_1 : boolean;
  signal phi_stmt_141_req_0 : boolean;
  signal phi_stmt_141_ack_0 : boolean;
  signal my_fetch4_99_143_buf_req_0 : boolean;
  signal my_fetch4_99_143_buf_ack_0 : boolean;
  signal my_fetch4_99_143_buf_req_1 : boolean;
  signal my_fetch4_99_143_buf_ack_1 : boolean;
  signal n_fetch_val4_492_144_buf_req_0 : boolean;
  signal n_fetch_val4_492_144_buf_ack_0 : boolean;
  signal n_fetch_val4_492_144_buf_req_1 : boolean;
  signal n_fetch_val4_492_144_buf_ack_1 : boolean;
  signal phi_stmt_145_req_1 : boolean;
  signal phi_stmt_145_req_0 : boolean;
  signal phi_stmt_145_ack_0 : boolean;
  signal n_row1_186_149_buf_req_0 : boolean;
  signal n_row1_186_149_buf_ack_0 : boolean;
  signal n_row1_186_149_buf_req_1 : boolean;
  signal n_row1_186_149_buf_ack_1 : boolean;
  signal phi_stmt_150_req_1 : boolean;
  signal phi_stmt_150_req_0 : boolean;
  signal phi_stmt_150_ack_0 : boolean;
  signal n_row2_194_154_buf_req_0 : boolean;
  signal n_row2_194_154_buf_ack_0 : boolean;
  signal n_row2_194_154_buf_req_1 : boolean;
  signal n_row2_194_154_buf_ack_1 : boolean;
  signal type_cast_227_inst_req_0 : boolean;
  signal type_cast_227_inst_ack_0 : boolean;
  signal type_cast_227_inst_req_1 : boolean;
  signal type_cast_227_inst_ack_1 : boolean;
  signal array_obj_ref_254_index_offset_req_0 : boolean;
  signal array_obj_ref_254_index_offset_ack_0 : boolean;
  signal array_obj_ref_254_index_offset_req_1 : boolean;
  signal array_obj_ref_254_index_offset_ack_1 : boolean;
  signal type_cast_371_inst_ack_1 : boolean;
  signal array_obj_ref_398_index_offset_req_0 : boolean;
  signal array_obj_ref_398_index_offset_ack_0 : boolean;
  signal array_obj_ref_398_index_offset_req_1 : boolean;
  signal array_obj_ref_398_index_offset_ack_1 : boolean;
  signal addr_of_399_final_reg_req_0 : boolean;
  signal addr_of_399_final_reg_ack_0 : boolean;
  signal addr_of_399_final_reg_req_1 : boolean;
  signal addr_of_399_final_reg_ack_1 : boolean;
  signal W_fn3_374_delayed_7_0_401_inst_req_0 : boolean;
  signal W_fn3_374_delayed_7_0_401_inst_ack_0 : boolean;
  signal W_fn3_374_delayed_7_0_401_inst_req_1 : boolean;
  signal W_fn3_374_delayed_7_0_401_inst_ack_1 : boolean;
  signal ptr_deref_407_load_0_req_0 : boolean;
  signal ptr_deref_407_load_0_ack_0 : boolean;
  signal ptr_deref_407_load_0_req_1 : boolean;
  signal ptr_deref_407_load_0_ack_1 : boolean;
  signal W_fn3_380_delayed_13_0_409_inst_req_0 : boolean;
  signal W_fn3_380_delayed_13_0_409_inst_ack_0 : boolean;
  signal W_fn3_380_delayed_13_0_409_inst_req_1 : boolean;
  signal W_fn3_380_delayed_13_0_409_inst_ack_1 : boolean;
  signal W_fetch_val3_382_delayed_13_0_412_inst_req_0 : boolean;
  signal W_fetch_val3_382_delayed_13_0_412_inst_ack_0 : boolean;
  signal W_fetch_val3_382_delayed_13_0_412_inst_req_1 : boolean;
  signal W_fetch_val3_382_delayed_13_0_412_inst_ack_1 : boolean;
  signal type_cast_443_inst_req_0 : boolean;
  signal type_cast_443_inst_ack_0 : boolean;
  signal type_cast_443_inst_req_1 : boolean;
  signal type_cast_443_inst_ack_1 : boolean;
  signal array_obj_ref_470_index_offset_req_0 : boolean;
  signal array_obj_ref_470_index_offset_ack_0 : boolean;
  signal array_obj_ref_470_index_offset_req_1 : boolean;
  signal array_obj_ref_470_index_offset_ack_1 : boolean;
  signal addr_of_471_final_reg_req_0 : boolean;
  signal addr_of_471_final_reg_ack_0 : boolean;
  signal addr_of_471_final_reg_req_1 : boolean;
  signal addr_of_471_final_reg_ack_1 : boolean;
  signal W_fn4_434_delayed_7_0_473_inst_req_0 : boolean;
  signal W_fn4_434_delayed_7_0_473_inst_ack_0 : boolean;
  signal W_fn4_434_delayed_7_0_473_inst_req_1 : boolean;
  signal W_fn4_434_delayed_7_0_473_inst_ack_1 : boolean;
  signal ptr_deref_479_load_0_req_0 : boolean;
  signal ptr_deref_479_load_0_ack_0 : boolean;
  signal ptr_deref_479_load_0_req_1 : boolean;
  signal ptr_deref_479_load_0_ack_1 : boolean;
  signal W_fn4_440_delayed_13_0_481_inst_req_0 : boolean;
  signal W_fn4_440_delayed_13_0_481_inst_ack_0 : boolean;
  signal W_fn4_440_delayed_13_0_481_inst_req_1 : boolean;
  signal W_fn4_440_delayed_13_0_481_inst_ack_1 : boolean;
  signal W_fetch_val4_442_delayed_13_0_484_inst_req_0 : boolean;
  signal W_fetch_val4_442_delayed_13_0_484_inst_ack_0 : boolean;
  signal W_fetch_val4_442_delayed_13_0_484_inst_req_1 : boolean;
  signal W_fetch_val4_442_delayed_13_0_484_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_494_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_494_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_494_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_494_inst_ack_1 : boolean;
  signal WPIPE_input_pipe2_498_inst_req_0 : boolean;
  signal WPIPE_input_pipe2_498_inst_ack_0 : boolean;
  signal WPIPE_input_pipe2_498_inst_req_1 : boolean;
  signal WPIPE_input_pipe2_498_inst_ack_1 : boolean;
  signal WPIPE_input_pipe3_502_inst_req_0 : boolean;
  signal WPIPE_input_pipe3_502_inst_ack_0 : boolean;
  signal WPIPE_input_pipe3_502_inst_req_1 : boolean;
  signal WPIPE_input_pipe3_502_inst_ack_1 : boolean;
  signal WPIPE_input_pipe4_506_inst_req_0 : boolean;
  signal WPIPE_input_pipe4_506_inst_ack_0 : boolean;
  signal WPIPE_input_pipe4_506_inst_req_1 : boolean;
  signal WPIPE_input_pipe4_506_inst_ack_1 : boolean;
  signal do_while_stmt_100_branch_ack_0 : boolean;
  signal do_while_stmt_100_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 48) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= row_in;
  row_in_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= ct;
  ct_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(tag_length + 47 downto 48) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 47 downto 48);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(377 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	19 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	17 
    -- CP-element group 0:  members (103) 
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_29/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/branch_block_stmt_29__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_complete/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_complete/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_complete/req
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_update_start_
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/word_0/cr
      -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_52_load_0_req_0); -- 
    cr_58_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_58_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_52_load_0_req_1); -- 
    req_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_75_index_offset_req_0); -- 
    req_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_61_index_offset_req_0); -- 
    req_94_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_94_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_61_index_offset_req_1); -- 
    req_109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_62_final_reg_req_1); -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_66_load_0_req_1); -- 
    req_190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_75_index_offset_req_1); -- 
    req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_76_final_reg_req_1); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_80_load_0_req_1); -- 
    req_281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_93_index_offset_req_0); -- 
    req_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_93_index_offset_req_1); -- 
    req_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_94_final_reg_req_1); -- 
    cr_346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_98_load_0_req_1); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	377 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_29/do_while_stmt_100__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_29/$exit
      -- CP-element group 1: 	 branch_block_stmt_29/branch_block_stmt_29__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(377);
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Sample/word_access_start/word_0/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_52_load_0_ack_0, ack => access_T_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	22 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/word_access_complete/word_0/ca
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/ptr_deref_52_Merge/$entry
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/ptr_deref_52_Merge/$exit
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/ptr_deref_52_Merge/merge_req
      -- CP-element group 3: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_52_Update/ptr_deref_52_Merge/merge_ack
      -- 
    ca_59_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_52_load_0_ack_1, ack => access_T_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	22 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_sample_complete
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Sample/ack
      -- 
    ack_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_index_offset_ack_0, ack => access_T_CP_0_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (11) 
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_root_address_calculated
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_offset_calculated
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_final_index_sum_regn_Update/ack
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_base_plus_offset/$entry
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_base_plus_offset/$exit
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_base_plus_offset/sum_rename_req
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_61_base_plus_offset/sum_rename_ack
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_request/$entry
      -- CP-element group 5: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_request/req
      -- 
    ack_95_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_61_index_offset_ack_1, ack => access_T_CP_0_elements(5)); -- 
    req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(5), ack => addr_of_62_final_reg_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_request/$exit
      -- CP-element group 6: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_request/ack
      -- 
    ack_105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_62_final_reg_ack_0, ack => access_T_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (24) 
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_62_complete/ack
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_root_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_address_resized
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_addr_resize/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_addr_resize/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_addr_resize/base_resize_req
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_addr_resize/base_resize_ack
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_plus_offset/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_plus_offset/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_plus_offset/sum_rename_req
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_base_plus_offset/sum_rename_ack
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_addrgen/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_addrgen/$exit
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_addrgen/root_register_req
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_word_addrgen/root_register_ack
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/word_0/rr
      -- 
    ack_110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_62_final_reg_ack_1, ack => access_T_CP_0_elements(7)); -- 
    rr_143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(7), ack => ptr_deref_66_load_0_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/$exit
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Sample/word_access_start/word_0/ra
      -- 
    ra_144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_load_0_ack_0, ack => access_T_CP_0_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	22 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/ptr_deref_66_Merge/$entry
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/ptr_deref_66_Merge/$exit
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/ptr_deref_66_Merge/merge_req
      -- CP-element group 9: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_66_Update/ptr_deref_66_Merge/merge_ack
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_load_0_ack_1, ack => access_T_CP_0_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	22 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_sample_complete
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Sample/ack
      -- 
    ack_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_75_index_offset_ack_0, ack => access_T_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (11) 
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_offset_calculated
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_final_index_sum_regn_Update/ack
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_base_plus_offset/$entry
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_base_plus_offset/$exit
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_base_plus_offset/sum_rename_req
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_75_base_plus_offset/sum_rename_ack
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_request/$entry
      -- CP-element group 11: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_request/req
      -- 
    ack_191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_75_index_offset_ack_1, ack => access_T_CP_0_elements(11)); -- 
    req_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(11), ack => addr_of_76_final_reg_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_request/$exit
      -- CP-element group 12: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_request/ack
      -- 
    ack_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_76_final_reg_ack_0, ack => access_T_CP_0_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (24) 
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_76_complete/ack
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_address_resized
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_addr_resize/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_addr_resize/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_addr_resize/base_resize_req
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_addr_resize/base_resize_ack
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_addrgen/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_addrgen/$exit
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_addrgen/root_register_req
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_word_addrgen/root_register_ack
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/word_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/word_0/rr
      -- 
    ack_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_76_final_reg_ack_1, ack => access_T_CP_0_elements(13)); -- 
    rr_239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(13), ack => ptr_deref_80_load_0_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/$exit
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Sample/word_access_start/word_0/ra
      -- 
    ra_240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_80_load_0_ack_0, ack => access_T_CP_0_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	22 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/word_access_complete/word_0/ca
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/ptr_deref_80_Merge/$entry
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/ptr_deref_80_Merge/$exit
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/ptr_deref_80_Merge/merge_req
      -- CP-element group 15: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_80_Update/ptr_deref_80_Merge/merge_ack
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_80_load_0_ack_1, ack => access_T_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_sample_complete
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Sample/ack
      -- 
    ack_282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_93_index_offset_ack_0, ack => access_T_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (11) 
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_root_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_offset_calculated
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_final_index_sum_regn_Update/ack
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_base_plus_offset/$entry
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_base_plus_offset/$exit
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/array_obj_ref_93_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_request/$entry
      -- CP-element group 17: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_request/req
      -- 
    ack_287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_93_index_offset_ack_1, ack => access_T_CP_0_elements(17)); -- 
    req_296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(17), ack => addr_of_94_final_reg_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_request/$exit
      -- CP-element group 18: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_request/ack
      -- 
    ack_297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_94_final_reg_ack_0, ack => access_T_CP_0_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	0 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (24) 
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/addr_of_94_complete/ack
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_root_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_address_resized
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_addr_resize/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_addr_resize/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_addr_resize/base_resize_req
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_addr_resize/base_resize_ack
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_plus_offset/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_plus_offset/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_base_plus_offset/sum_rename_ack
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_addrgen/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_addrgen/$exit
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_addrgen/root_register_req
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_word_addrgen/root_register_ack
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/word_0/rr
      -- 
    ack_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_94_final_reg_ack_1, ack => access_T_CP_0_elements(19)); -- 
    rr_335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(19), ack => ptr_deref_98_load_0_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Sample/word_access_start/word_0/ra
      -- 
    ra_336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_98_load_0_ack_0, ack => access_T_CP_0_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/ptr_deref_98_Merge/$entry
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/ptr_deref_98_Merge/$exit
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/ptr_deref_98_Merge/merge_req
      -- CP-element group 21: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/ptr_deref_98_Update/ptr_deref_98_Merge/merge_ack
      -- 
    ca_347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_98_load_0_ack_1, ack => access_T_CP_0_elements(21)); -- 
    -- CP-element group 22:  join  transition  place  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: 	3 
    -- CP-element group 22: 	4 
    -- CP-element group 22: 	9 
    -- CP-element group 22: 	10 
    -- CP-element group 22: 	15 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99__exit__
      -- CP-element group 22: 	 branch_block_stmt_29/do_while_stmt_100__entry__
      -- CP-element group 22: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_99/$exit
      -- 
    access_T_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(21) & access_T_CP_0_elements(3) & access_T_CP_0_elements(4) & access_T_CP_0_elements(9) & access_T_CP_0_elements(10) & access_T_CP_0_elements(15) & access_T_CP_0_elements(16);
      gj_access_T_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  place  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	29 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_29/do_while_stmt_100/$entry
      -- CP-element group 23: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100__entry__
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(22);
    -- CP-element group 24:  merge  place  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	377 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100__exit__
      -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  merge  place  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_29/do_while_stmt_100/loop_back
      -- 
    -- Element group access_T_CP_0_elements(25) is bound as output of CP function.
    -- CP-element group 26:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	375 
    -- CP-element group 26: 	376 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_100/condition_done
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_100/loop_exit/$entry
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_100/loop_taken/$entry
      -- 
    access_T_CP_0_elements(26) <= access_T_CP_0_elements(31);
    -- CP-element group 27:  branch  place  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	374 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_29/do_while_stmt_100/loop_body_done
      -- 
    access_T_CP_0_elements(27) <= access_T_CP_0_elements(374);
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	80 
    -- CP-element group 28: 	101 
    -- CP-element group 28: 	122 
    -- CP-element group 28: 	42 
    -- CP-element group 28: 	61 
    -- CP-element group 28: 	141 
    -- CP-element group 28: 	160 
    -- CP-element group 28: 	179 
    -- CP-element group 28: 	198 
    -- CP-element group 28: 	217 
    -- CP-element group 28: 	236 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(28) <= access_T_CP_0_elements(25);
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	103 
    -- CP-element group 29: 	124 
    -- CP-element group 29: 	44 
    -- CP-element group 29: 	63 
    -- CP-element group 29: 	82 
    -- CP-element group 29: 	143 
    -- CP-element group 29: 	162 
    -- CP-element group 29: 	181 
    -- CP-element group 29: 	200 
    -- CP-element group 29: 	219 
    -- CP-element group 29: 	238 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(29) <= access_T_CP_0_elements(23);
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	76 
    -- CP-element group 30: 	77 
    -- CP-element group 30: 	95 
    -- CP-element group 30: 	96 
    -- CP-element group 30: 	116 
    -- CP-element group 30: 	117 
    -- CP-element group 30: 	135 
    -- CP-element group 30: 	136 
    -- CP-element group 30: 	56 
    -- CP-element group 30: 	36 
    -- CP-element group 30: 	37 
    -- CP-element group 30: 	55 
    -- CP-element group 30: 	154 
    -- CP-element group 30: 	155 
    -- CP-element group 30: 	173 
    -- CP-element group 30: 	174 
    -- CP-element group 30: 	192 
    -- CP-element group 30: 	193 
    -- CP-element group 30: 	211 
    -- CP-element group 30: 	212 
    -- CP-element group 30: 	230 
    -- CP-element group 30: 	231 
    -- CP-element group 30: 	249 
    -- CP-element group 30: 	254 
    -- CP-element group 30: 	256 
    -- CP-element group 30: 	277 
    -- CP-element group 30: 	282 
    -- CP-element group 30: 	284 
    -- CP-element group 30: 	305 
    -- CP-element group 30: 	310 
    -- CP-element group 30: 	312 
    -- CP-element group 30: 	333 
    -- CP-element group 30: 	338 
    -- CP-element group 30: 	340 
    -- CP-element group 30: 	373 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/$entry
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	121 
    -- CP-element group 31: 	35 
    -- CP-element group 31: 	216 
    -- CP-element group 31: 	373 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	26 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/condition_evaluated
      -- 
    condition_evaluated_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(31), ack => do_while_stmt_100_branch_req_0); -- 
    access_T_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(121) & access_T_CP_0_elements(35) & access_T_CP_0_elements(216) & access_T_CP_0_elements(373);
      gj_access_T_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	76 
    -- CP-element group 32: 	95 
    -- CP-element group 32: 	116 
    -- CP-element group 32: 	135 
    -- CP-element group 32: 	36 
    -- CP-element group 32: 	55 
    -- CP-element group 32: 	154 
    -- CP-element group 32: 	173 
    -- CP-element group 32: 	192 
    -- CP-element group 32: 	211 
    -- CP-element group 32: 	230 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	35 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	97 
    -- CP-element group 32: 	118 
    -- CP-element group 32: 	137 
    -- CP-element group 32: 	38 
    -- CP-element group 32: 	57 
    -- CP-element group 32: 	156 
    -- CP-element group 32: 	175 
    -- CP-element group 32: 	194 
    -- CP-element group 32: 	213 
    -- CP-element group 32: 	232 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/aggregated_phi_sample_req
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_sample_start__ps
      -- 
    access_T_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= access_T_CP_0_elements(76) & access_T_CP_0_elements(95) & access_T_CP_0_elements(116) & access_T_CP_0_elements(135) & access_T_CP_0_elements(36) & access_T_CP_0_elements(55) & access_T_CP_0_elements(154) & access_T_CP_0_elements(173) & access_T_CP_0_elements(192) & access_T_CP_0_elements(211) & access_T_CP_0_elements(230) & access_T_CP_0_elements(35);
      gj_access_T_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	98 
    -- CP-element group 33: 	119 
    -- CP-element group 33: 	138 
    -- CP-element group 33: 	39 
    -- CP-element group 33: 	58 
    -- CP-element group 33: 	157 
    -- CP-element group 33: 	176 
    -- CP-element group 33: 	195 
    -- CP-element group 33: 	214 
    -- CP-element group 33: 	233 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	250 
    -- CP-element group 33: 	266 
    -- CP-element group 33: 	270 
    -- CP-element group 33: 	274 
    -- CP-element group 33: 	278 
    -- CP-element group 33: 	294 
    -- CP-element group 33: 	298 
    -- CP-element group 33: 	302 
    -- CP-element group 33: 	306 
    -- CP-element group 33: 	322 
    -- CP-element group 33: 	326 
    -- CP-element group 33: 	330 
    -- CP-element group 33: 	334 
    -- CP-element group 33: 	350 
    -- CP-element group 33: 	354 
    -- CP-element group 33: 	358 
    -- CP-element group 33: 	374 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	76 
    -- CP-element group 33: 	95 
    -- CP-element group 33: 	116 
    -- CP-element group 33: 	135 
    -- CP-element group 33: 	36 
    -- CP-element group 33: 	55 
    -- CP-element group 33: 	154 
    -- CP-element group 33: 	173 
    -- CP-element group 33: 	192 
    -- CP-element group 33: 	211 
    -- CP-element group 33: 	230 
    -- CP-element group 33:  members (12) 
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/aggregated_phi_sample_ack
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_sample_completed_
      -- 
    access_T_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(78) & access_T_CP_0_elements(98) & access_T_CP_0_elements(119) & access_T_CP_0_elements(138) & access_T_CP_0_elements(39) & access_T_CP_0_elements(58) & access_T_CP_0_elements(157) & access_T_CP_0_elements(176) & access_T_CP_0_elements(195) & access_T_CP_0_elements(214) & access_T_CP_0_elements(233);
      gj_access_T_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	77 
    -- CP-element group 34: 	96 
    -- CP-element group 34: 	117 
    -- CP-element group 34: 	136 
    -- CP-element group 34: 	56 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	155 
    -- CP-element group 34: 	174 
    -- CP-element group 34: 	193 
    -- CP-element group 34: 	212 
    -- CP-element group 34: 	231 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	99 
    -- CP-element group 34: 	120 
    -- CP-element group 34: 	139 
    -- CP-element group 34: 	59 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	158 
    -- CP-element group 34: 	177 
    -- CP-element group 34: 	196 
    -- CP-element group 34: 	215 
    -- CP-element group 34: 	234 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/aggregated_phi_update_req
      -- CP-element group 34: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_update_start__ps
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(77) & access_T_CP_0_elements(96) & access_T_CP_0_elements(117) & access_T_CP_0_elements(136) & access_T_CP_0_elements(56) & access_T_CP_0_elements(37) & access_T_CP_0_elements(155) & access_T_CP_0_elements(174) & access_T_CP_0_elements(193) & access_T_CP_0_elements(212) & access_T_CP_0_elements(231);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	79 
    -- CP-element group 35: 	100 
    -- CP-element group 35: 	121 
    -- CP-element group 35: 	60 
    -- CP-element group 35: 	41 
    -- CP-element group 35: 	140 
    -- CP-element group 35: 	159 
    -- CP-element group 35: 	178 
    -- CP-element group 35: 	197 
    -- CP-element group 35: 	216 
    -- CP-element group 35: 	235 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	31 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	32 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(79) & access_T_CP_0_elements(100) & access_T_CP_0_elements(121) & access_T_CP_0_elements(60) & access_T_CP_0_elements(41) & access_T_CP_0_elements(140) & access_T_CP_0_elements(159) & access_T_CP_0_elements(178) & access_T_CP_0_elements(197) & access_T_CP_0_elements(216) & access_T_CP_0_elements(235);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	30 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	252 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	32 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_sample_start_
      -- 
    access_T_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(252);
      gj_access_T_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	30 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	41 
    -- CP-element group 37: 	257 
    -- CP-element group 37: 	263 
    -- CP-element group 37: 	271 
    -- CP-element group 37: 	362 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	34 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_update_start_
      -- 
    access_T_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(41) & access_T_CP_0_elements(257) & access_T_CP_0_elements(263) & access_T_CP_0_elements(271) & access_T_CP_0_elements(362);
      gj_access_T_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_sample_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(32);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	33 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_update_start__ps
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(34);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	35 
    -- CP-element group 41: 	255 
    -- CP-element group 41: 	261 
    -- CP-element group 41: 	269 
    -- CP-element group 41: 	361 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	37 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	28 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_loopback_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(28);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_loopback_sample_req_ps
      -- 
    phi_stmt_102_loopback_sample_req_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_102_loopback_sample_req_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_102_req_1); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	29 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_entry_trigger
      -- 
    access_T_CP_0_elements(44) <= access_T_CP_0_elements(29);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_entry_sample_req
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_entry_sample_req_ps
      -- 
    phi_stmt_102_entry_sample_req_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_102_entry_sample_req_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(45), ack => phi_stmt_102_req_0); -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_102_phi_mux_ack_ps
      -- 
    phi_stmt_102_phi_mux_ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_102_ack_0, ack => access_T_CP_0_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_update_start_
      -- 
    -- Element group access_T_CP_0_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_update_completed__ps
      -- 
    access_T_CP_0_elements(49) <= access_T_CP_0_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_105_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(48), ack => access_T_CP_0_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_sample_start__ps
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Sample/req
      -- 
    req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(51), ack => n_address1_236_106_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_update_start__ps
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_update_start_
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Update/req
      -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(52), ack => n_address1_236_106_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Sample/ack
      -- 
    ack_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_236_106_buf_ack_0, ack => access_T_CP_0_elements(53)); -- 
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address1_106_Update/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_236_106_buf_ack_1, ack => access_T_CP_0_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	30 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	33 
    -- CP-element group 55: 	280 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	32 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_sample_start_
      -- 
    access_T_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(280);
      gj_access_T_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	30 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	285 
    -- CP-element group 56: 	291 
    -- CP-element group 56: 	299 
    -- CP-element group 56: 	365 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	34 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_update_start_
      -- 
    access_T_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(60) & access_T_CP_0_elements(285) & access_T_CP_0_elements(291) & access_T_CP_0_elements(299) & access_T_CP_0_elements(365);
      gj_access_T_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	32 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_sample_start__ps
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(32);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	33 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	34 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_update_start__ps
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(34);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	35 
    -- CP-element group 60: 	283 
    -- CP-element group 60: 	289 
    -- CP-element group 60: 	297 
    -- CP-element group 60: 	364 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	56 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	28 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_loopback_trigger
      -- 
    access_T_CP_0_elements(61) <= access_T_CP_0_elements(28);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_loopback_sample_req_ps
      -- 
    phi_stmt_107_loopback_sample_req_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_107_loopback_sample_req_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => phi_stmt_107_req_1); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	29 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_entry_trigger
      -- 
    access_T_CP_0_elements(63) <= access_T_CP_0_elements(29);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_entry_sample_req_ps
      -- 
    phi_stmt_107_entry_sample_req_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_107_entry_sample_req_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => phi_stmt_107_req_0); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_107_phi_mux_ack_ps
      -- 
    phi_stmt_107_phi_mux_ack_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_107_ack_0, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Sample/rr
      -- 
    rr_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(68), ack => type_cast_110_inst_req_0); -- 
    access_T_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(66) & access_T_CP_0_elements(70);
      gj_access_T_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_update_start_
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Update/cr
      -- 
    cr_450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(69), ack => type_cast_110_inst_req_1); -- 
    access_T_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(67) & access_T_CP_0_elements(71);
      gj_access_T_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Sample/ra
      -- 
    ra_446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_0, ack => access_T_CP_0_elements(70)); -- 
    -- CP-element group 71:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_110_Update/ca
      -- 
    ca_451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_1, ack => access_T_CP_0_elements(71)); -- 
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_sample_start__ps
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Sample/req
      -- 
    req_463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(72), ack => n_address2_308_111_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_update_start__ps
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_update_start_
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Update/req
      -- 
    req_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(73), ack => n_address2_308_111_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_sample_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Sample/ack
      -- 
    ack_464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_308_111_buf_ack_0, ack => access_T_CP_0_elements(74)); -- 
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address2_111_Update/ack
      -- 
    ack_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_308_111_buf_ack_1, ack => access_T_CP_0_elements(75)); -- 
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	30 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	33 
    -- CP-element group 76: 	308 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	32 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_sample_start_
      -- 
    access_T_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(308);
      gj_access_T_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	30 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	313 
    -- CP-element group 77: 	319 
    -- CP-element group 77: 	327 
    -- CP-element group 77: 	368 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	34 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_update_start_
      -- 
    access_T_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(79) & access_T_CP_0_elements(313) & access_T_CP_0_elements(319) & access_T_CP_0_elements(327) & access_T_CP_0_elements(368);
      gj_access_T_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	33 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(78) is bound as output of CP function.
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	35 
    -- CP-element group 79: 	311 
    -- CP-element group 79: 	317 
    -- CP-element group 79: 	325 
    -- CP-element group 79: 	367 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	28 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_loopback_trigger
      -- 
    access_T_CP_0_elements(80) <= access_T_CP_0_elements(28);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_loopback_sample_req
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_loopback_sample_req_ps
      -- 
    phi_stmt_112_loopback_sample_req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_112_loopback_sample_req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(81), ack => phi_stmt_112_req_1); -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	29 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_entry_trigger
      -- 
    access_T_CP_0_elements(82) <= access_T_CP_0_elements(29);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_entry_sample_req
      -- CP-element group 83: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_entry_sample_req_ps
      -- 
    phi_stmt_112_entry_sample_req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_112_entry_sample_req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => phi_stmt_112_req_0); -- 
    -- Element group access_T_CP_0_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_phi_mux_ack
      -- CP-element group 84: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_112_phi_mux_ack_ps
      -- 
    phi_stmt_112_phi_mux_ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_112_ack_0, ack => access_T_CP_0_elements(84)); -- 
    -- CP-element group 85:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Sample/rr
      -- 
    rr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(87), ack => type_cast_115_inst_req_0); -- 
    access_T_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(85) & access_T_CP_0_elements(89);
      gj_access_T_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_update_start_
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Update/cr
      -- 
    cr_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(88), ack => type_cast_115_inst_req_1); -- 
    access_T_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(86) & access_T_CP_0_elements(90);
      gj_access_T_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Sample/ra
      -- 
    ra_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_0, ack => access_T_CP_0_elements(89)); -- 
    -- CP-element group 90:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_115_Update/ca
      -- 
    ca_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_1, ack => access_T_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_sample_start__ps
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Sample/req
      -- 
    req_517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(91), ack => n_address3_380_116_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(91) is bound as output of CP function.
    -- CP-element group 92:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_update_start__ps
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_update_start_
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Update/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(92), ack => n_address3_380_116_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_sample_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Sample/ack
      -- 
    ack_518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_380_116_buf_ack_0, ack => access_T_CP_0_elements(93)); -- 
    -- CP-element group 94:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_update_completed__ps
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address3_116_Update/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_380_116_buf_ack_1, ack => access_T_CP_0_elements(94)); -- 
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	30 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	33 
    -- CP-element group 95: 	336 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	32 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_sample_start_
      -- 
    access_T_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(336);
      gj_access_T_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	30 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	100 
    -- CP-element group 96: 	341 
    -- CP-element group 96: 	347 
    -- CP-element group 96: 	355 
    -- CP-element group 96: 	371 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	34 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_update_start_
      -- 
    access_T_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(100) & access_T_CP_0_elements(341) & access_T_CP_0_elements(347) & access_T_CP_0_elements(355) & access_T_CP_0_elements(371);
      gj_access_T_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	32 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_sample_start__ps
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(32);
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	33 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	34 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_update_start__ps
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(34);
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	35 
    -- CP-element group 100: 	339 
    -- CP-element group 100: 	345 
    -- CP-element group 100: 	353 
    -- CP-element group 100: 	370 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	96 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	28 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_loopback_trigger
      -- 
    access_T_CP_0_elements(101) <= access_T_CP_0_elements(28);
    -- CP-element group 102:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_loopback_sample_req
      -- CP-element group 102: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_loopback_sample_req_ps
      -- 
    phi_stmt_117_loopback_sample_req_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_117_loopback_sample_req_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(102), ack => phi_stmt_117_req_1); -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	29 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_entry_trigger
      -- 
    access_T_CP_0_elements(103) <= access_T_CP_0_elements(29);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_entry_sample_req
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_entry_sample_req_ps
      -- 
    phi_stmt_117_entry_sample_req_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_117_entry_sample_req_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(104), ack => phi_stmt_117_req_0); -- 
    -- Element group access_T_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_phi_mux_ack
      -- CP-element group 105: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_117_phi_mux_ack_ps
      -- 
    phi_stmt_117_phi_mux_ack_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_117_ack_0, ack => access_T_CP_0_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Sample/rr
      -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(108), ack => type_cast_122_inst_req_0); -- 
    access_T_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(106) & access_T_CP_0_elements(110);
      gj_access_T_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_update_start_
      -- CP-element group 109: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Update/cr
      -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(109), ack => type_cast_122_inst_req_1); -- 
    access_T_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(107) & access_T_CP_0_elements(111);
      gj_access_T_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (4) 
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_sample_completed__ps
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Sample/ra
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_122_inst_ack_0, ack => access_T_CP_0_elements(110)); -- 
    -- CP-element group 111:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_update_completed__ps
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_122_Update/ca
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_122_inst_ack_1, ack => access_T_CP_0_elements(111)); -- 
    -- CP-element group 112:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_sample_start__ps
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Sample/req
      -- 
    req_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(112), ack => n_address4_452_123_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_update_start__ps
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_update_start_
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Update/req
      -- 
    req_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(113), ack => n_address4_452_123_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Sample/ack
      -- 
    ack_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address4_452_123_buf_ack_0, ack => access_T_CP_0_elements(114)); -- 
    -- CP-element group 115:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_update_completed__ps
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_address4_123_Update/ack
      -- 
    ack_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address4_452_123_buf_ack_1, ack => access_T_CP_0_elements(115)); -- 
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	30 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	33 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	32 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_sample_start_
      -- 
    access_T_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33);
      gj_access_T_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	30 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: 	257 
    -- CP-element group 117: 	263 
    -- CP-element group 117: 	271 
    -- CP-element group 117: 	285 
    -- CP-element group 117: 	291 
    -- CP-element group 117: 	299 
    -- CP-element group 117: 	313 
    -- CP-element group 117: 	319 
    -- CP-element group 117: 	327 
    -- CP-element group 117: 	341 
    -- CP-element group 117: 	347 
    -- CP-element group 117: 	355 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	34 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_update_start_
      -- 
    access_T_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 1,6 => 0,7 => 0,8 => 1,9 => 0,10 => 0,11 => 1,12 => 0,13 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(121) & access_T_CP_0_elements(257) & access_T_CP_0_elements(263) & access_T_CP_0_elements(271) & access_T_CP_0_elements(285) & access_T_CP_0_elements(291) & access_T_CP_0_elements(299) & access_T_CP_0_elements(313) & access_T_CP_0_elements(319) & access_T_CP_0_elements(327) & access_T_CP_0_elements(341) & access_T_CP_0_elements(347) & access_T_CP_0_elements(355);
      gj_access_T_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	32 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_sample_start__ps
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(32);
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	33 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	34 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_update_start__ps
      -- 
    access_T_CP_0_elements(120) <= access_T_CP_0_elements(34);
    -- CP-element group 121:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	35 
    -- CP-element group 121: 	31 
    -- CP-element group 121: 	255 
    -- CP-element group 121: 	261 
    -- CP-element group 121: 	269 
    -- CP-element group 121: 	283 
    -- CP-element group 121: 	289 
    -- CP-element group 121: 	297 
    -- CP-element group 121: 	311 
    -- CP-element group 121: 	317 
    -- CP-element group 121: 	325 
    -- CP-element group 121: 	339 
    -- CP-element group 121: 	345 
    -- CP-element group 121: 	353 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	117 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	28 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_loopback_trigger
      -- 
    access_T_CP_0_elements(122) <= access_T_CP_0_elements(28);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_loopback_sample_req
      -- CP-element group 123: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_loopback_sample_req_ps
      -- 
    phi_stmt_124_loopback_sample_req_588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_124_loopback_sample_req_588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(123), ack => phi_stmt_124_req_1); -- 
    -- Element group access_T_CP_0_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	29 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_entry_trigger
      -- 
    access_T_CP_0_elements(124) <= access_T_CP_0_elements(29);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_entry_sample_req
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_entry_sample_req_ps
      -- 
    phi_stmt_124_entry_sample_req_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_124_entry_sample_req_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => phi_stmt_124_req_0); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_phi_mux_ack
      -- CP-element group 126: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_124_phi_mux_ack_ps
      -- 
    phi_stmt_124_phi_mux_ack_594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_124_ack_0, ack => access_T_CP_0_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_sample_start__ps
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_update_start__ps
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_update_start_
      -- 
    -- Element group access_T_CP_0_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_update_completed__ps
      -- 
    access_T_CP_0_elements(129) <= access_T_CP_0_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_127_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(128), ack => access_T_CP_0_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_sample_start__ps
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Sample/req
      -- 
    req_615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(131), ack => n_mycounter_168_128_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_update_start__ps
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_update_start_
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Update/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(132), ack => n_mycounter_168_128_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Sample/ack
      -- 
    ack_616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter_168_128_buf_ack_0, ack => access_T_CP_0_elements(133)); -- 
    -- CP-element group 134:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_mycounter_128_Update/ack
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter_168_128_buf_ack_1, ack => access_T_CP_0_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	30 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	33 
    -- CP-element group 135: 	268 
    -- CP-element group 135: 	272 
    -- CP-element group 135: 	276 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	32 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_sample_start_
      -- 
    access_T_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(268) & access_T_CP_0_elements(272) & access_T_CP_0_elements(276);
      gj_access_T_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	30 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	140 
    -- CP-element group 136: 	275 
    -- CP-element group 136: 	362 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	34 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_update_start_
      -- 
    access_T_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(140) & access_T_CP_0_elements(275) & access_T_CP_0_elements(362);
      gj_access_T_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	32 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_sample_start__ps
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(32);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	33 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	34 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_update_start__ps
      -- 
    access_T_CP_0_elements(139) <= access_T_CP_0_elements(34);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	35 
    -- CP-element group 140: 	273 
    -- CP-element group 140: 	361 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	136 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	28 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_loopback_trigger
      -- 
    access_T_CP_0_elements(141) <= access_T_CP_0_elements(28);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_loopback_sample_req_ps
      -- 
    phi_stmt_129_loopback_sample_req_632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_129_loopback_sample_req_632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(142), ack => phi_stmt_129_req_1); -- 
    -- Element group access_T_CP_0_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	29 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_entry_trigger
      -- 
    access_T_CP_0_elements(143) <= access_T_CP_0_elements(29);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_entry_sample_req_ps
      -- 
    phi_stmt_129_entry_sample_req_635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_129_entry_sample_req_635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(144), ack => phi_stmt_129_req_0); -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_129_phi_mux_ack_ps
      -- 
    phi_stmt_129_phi_mux_ack_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_129_ack_0, ack => access_T_CP_0_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Sample/req
      -- 
    req_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(146), ack => my_fetch1_53_131_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_update_start_
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Update/req
      -- 
    req_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(147), ack => my_fetch1_53_131_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (4) 
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_sample_completed__ps
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Sample/ack
      -- 
    ack_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch1_53_131_buf_ack_0, ack => access_T_CP_0_elements(148)); -- 
    -- CP-element group 149:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (4) 
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_update_completed__ps
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch1_131_Update/ack
      -- 
    ack_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch1_53_131_buf_ack_1, ack => access_T_CP_0_elements(149)); -- 
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_sample_start_
      -- 
    req_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => n_fetch_val1_276_132_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Update/req
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_update_start_
      -- 
    req_674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(151), ack => n_fetch_val1_276_132_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_sample_completed_
      -- 
    ack_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val1_276_132_buf_ack_0, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val1_132_update_completed__ps
      -- 
    ack_675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val1_276_132_buf_ack_1, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  join  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	30 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	33 
    -- CP-element group 154: 	296 
    -- CP-element group 154: 	300 
    -- CP-element group 154: 	304 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	32 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_sample_start_
      -- 
    access_T_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(296) & access_T_CP_0_elements(300) & access_T_CP_0_elements(304);
      gj_access_T_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	30 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	159 
    -- CP-element group 155: 	303 
    -- CP-element group 155: 	365 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	34 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_update_start_
      -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(159) & access_T_CP_0_elements(303) & access_T_CP_0_elements(365);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	32 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_sample_start__ps
      -- 
    access_T_CP_0_elements(156) <= access_T_CP_0_elements(32);
    -- CP-element group 157:  join  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	33 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(157) is bound as output of CP function.
    -- CP-element group 158:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	34 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_update_start__ps
      -- 
    access_T_CP_0_elements(158) <= access_T_CP_0_elements(34);
    -- CP-element group 159:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	35 
    -- CP-element group 159: 	301 
    -- CP-element group 159: 	364 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	155 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(159) is bound as output of CP function.
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	28 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_loopback_trigger
      -- 
    access_T_CP_0_elements(160) <= access_T_CP_0_elements(28);
    -- CP-element group 161:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (2) 
      -- CP-element group 161: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_loopback_sample_req
      -- CP-element group 161: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_loopback_sample_req_ps
      -- 
    phi_stmt_133_loopback_sample_req_686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_loopback_sample_req_686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(161), ack => phi_stmt_133_req_1); -- 
    -- Element group access_T_CP_0_elements(161) is bound as output of CP function.
    -- CP-element group 162:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	29 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_entry_trigger
      -- 
    access_T_CP_0_elements(162) <= access_T_CP_0_elements(29);
    -- CP-element group 163:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_entry_sample_req
      -- CP-element group 163: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_entry_sample_req_ps
      -- 
    phi_stmt_133_entry_sample_req_689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_133_entry_sample_req_689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => phi_stmt_133_req_0); -- 
    -- Element group access_T_CP_0_elements(163) is bound as output of CP function.
    -- CP-element group 164:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_phi_mux_ack
      -- CP-element group 164: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_133_phi_mux_ack_ps
      -- 
    phi_stmt_133_phi_mux_ack_692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_133_ack_0, ack => access_T_CP_0_elements(164)); -- 
    -- CP-element group 165:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (4) 
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_sample_start__ps
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Sample/req
      -- 
    req_705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(165), ack => my_fetch2_67_135_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(165) is bound as output of CP function.
    -- CP-element group 166:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (4) 
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_update_start__ps
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_update_start_
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Update/req
      -- 
    req_710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(166), ack => my_fetch2_67_135_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(166) is bound as output of CP function.
    -- CP-element group 167:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (4) 
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_sample_completed__ps
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Sample/ack
      -- 
    ack_706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch2_67_135_buf_ack_0, ack => access_T_CP_0_elements(167)); -- 
    -- CP-element group 168:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (4) 
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_update_completed__ps
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch2_135_Update/ack
      -- 
    ack_711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch2_67_135_buf_ack_1, ack => access_T_CP_0_elements(168)); -- 
    -- CP-element group 169:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (4) 
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_sample_start__ps
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Sample/req
      -- 
    req_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(169), ack => n_fetch_val2_348_136_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(169) is bound as output of CP function.
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_update_start__ps
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_update_start_
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Update/req
      -- 
    req_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(170), ack => n_fetch_val2_348_136_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (4) 
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_sample_completed__ps
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Sample/ack
      -- 
    ack_724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val2_348_136_buf_ack_0, ack => access_T_CP_0_elements(171)); -- 
    -- CP-element group 172:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (4) 
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_update_completed__ps
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val2_136_Update/ack
      -- 
    ack_729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val2_348_136_buf_ack_1, ack => access_T_CP_0_elements(172)); -- 
    -- CP-element group 173:  join  transition  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	30 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	33 
    -- CP-element group 173: 	324 
    -- CP-element group 173: 	328 
    -- CP-element group 173: 	332 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	32 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_sample_start_
      -- 
    access_T_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(324) & access_T_CP_0_elements(328) & access_T_CP_0_elements(332);
      gj_access_T_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	30 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	178 
    -- CP-element group 174: 	331 
    -- CP-element group 174: 	368 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	34 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_update_start_
      -- 
    access_T_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(178) & access_T_CP_0_elements(331) & access_T_CP_0_elements(368);
      gj_access_T_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	32 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_sample_start__ps
      -- 
    access_T_CP_0_elements(175) <= access_T_CP_0_elements(32);
    -- CP-element group 176:  join  transition  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	33 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(176) is bound as output of CP function.
    -- CP-element group 177:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	34 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_update_start__ps
      -- 
    access_T_CP_0_elements(177) <= access_T_CP_0_elements(34);
    -- CP-element group 178:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	35 
    -- CP-element group 178: 	329 
    -- CP-element group 178: 	367 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	174 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(178) is bound as output of CP function.
    -- CP-element group 179:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	28 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_loopback_trigger
      -- 
    access_T_CP_0_elements(179) <= access_T_CP_0_elements(28);
    -- CP-element group 180:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_loopback_sample_req
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_loopback_sample_req_ps
      -- 
    phi_stmt_137_loopback_sample_req_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_137_loopback_sample_req_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => phi_stmt_137_req_1); -- 
    -- Element group access_T_CP_0_elements(180) is bound as output of CP function.
    -- CP-element group 181:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	29 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_entry_trigger
      -- 
    access_T_CP_0_elements(181) <= access_T_CP_0_elements(29);
    -- CP-element group 182:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_entry_sample_req
      -- CP-element group 182: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_entry_sample_req_ps
      -- 
    phi_stmt_137_entry_sample_req_743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_137_entry_sample_req_743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => phi_stmt_137_req_0); -- 
    -- Element group access_T_CP_0_elements(182) is bound as output of CP function.
    -- CP-element group 183:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_phi_mux_ack
      -- CP-element group 183: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_137_phi_mux_ack_ps
      -- 
    phi_stmt_137_phi_mux_ack_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_137_ack_0, ack => access_T_CP_0_elements(183)); -- 
    -- CP-element group 184:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (4) 
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_sample_start__ps
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Sample/req
      -- 
    req_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(184), ack => my_fetch3_81_139_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(184) is bound as output of CP function.
    -- CP-element group 185:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (4) 
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_update_start__ps
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_update_start_
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Update/req
      -- 
    req_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(185), ack => my_fetch3_81_139_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(185) is bound as output of CP function.
    -- CP-element group 186:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (4) 
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_sample_completed__ps
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Sample/ack
      -- 
    ack_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch3_81_139_buf_ack_0, ack => access_T_CP_0_elements(186)); -- 
    -- CP-element group 187:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (4) 
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_update_completed__ps
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch3_139_Update/ack
      -- 
    ack_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch3_81_139_buf_ack_1, ack => access_T_CP_0_elements(187)); -- 
    -- CP-element group 188:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (4) 
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_sample_start__ps
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Sample/req
      -- 
    req_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(188), ack => n_fetch_val3_420_140_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(188) is bound as output of CP function.
    -- CP-element group 189:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (4) 
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_update_start__ps
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_update_start_
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Update/req
      -- 
    req_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => n_fetch_val3_420_140_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(189) is bound as output of CP function.
    -- CP-element group 190:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (4) 
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_sample_completed__ps
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Sample/ack
      -- 
    ack_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val3_420_140_buf_ack_0, ack => access_T_CP_0_elements(190)); -- 
    -- CP-element group 191:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (4) 
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_update_completed__ps
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val3_140_Update/ack
      -- 
    ack_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val3_420_140_buf_ack_1, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  join  transition  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	30 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	33 
    -- CP-element group 192: 	352 
    -- CP-element group 192: 	356 
    -- CP-element group 192: 	360 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	32 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_sample_start_
      -- 
    access_T_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33) & access_T_CP_0_elements(352) & access_T_CP_0_elements(356) & access_T_CP_0_elements(360);
      gj_access_T_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	30 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	197 
    -- CP-element group 193: 	359 
    -- CP-element group 193: 	371 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	34 
    -- CP-element group 193:  members (1) 
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_update_start_
      -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(197) & access_T_CP_0_elements(359) & access_T_CP_0_elements(371);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	32 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (1) 
      -- CP-element group 194: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_sample_start__ps
      -- 
    access_T_CP_0_elements(194) <= access_T_CP_0_elements(32);
    -- CP-element group 195:  join  transition  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	33 
    -- CP-element group 195:  members (1) 
      -- CP-element group 195: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(195) is bound as output of CP function.
    -- CP-element group 196:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	34 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_update_start__ps
      -- 
    access_T_CP_0_elements(196) <= access_T_CP_0_elements(34);
    -- CP-element group 197:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	35 
    -- CP-element group 197: 	357 
    -- CP-element group 197: 	370 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	193 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(197) is bound as output of CP function.
    -- CP-element group 198:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	28 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_loopback_trigger
      -- 
    access_T_CP_0_elements(198) <= access_T_CP_0_elements(28);
    -- CP-element group 199:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_loopback_sample_req
      -- CP-element group 199: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_loopback_sample_req_ps
      -- 
    phi_stmt_141_loopback_sample_req_794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_141_loopback_sample_req_794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(199), ack => phi_stmt_141_req_1); -- 
    -- Element group access_T_CP_0_elements(199) is bound as output of CP function.
    -- CP-element group 200:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	29 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_entry_trigger
      -- 
    access_T_CP_0_elements(200) <= access_T_CP_0_elements(29);
    -- CP-element group 201:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (2) 
      -- CP-element group 201: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_entry_sample_req
      -- CP-element group 201: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_entry_sample_req_ps
      -- 
    phi_stmt_141_entry_sample_req_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_141_entry_sample_req_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => phi_stmt_141_req_0); -- 
    -- Element group access_T_CP_0_elements(201) is bound as output of CP function.
    -- CP-element group 202:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (2) 
      -- CP-element group 202: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_phi_mux_ack
      -- CP-element group 202: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_141_phi_mux_ack_ps
      -- 
    phi_stmt_141_phi_mux_ack_800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_141_ack_0, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (4) 
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_sample_start__ps
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Sample/req
      -- 
    req_813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(203), ack => my_fetch4_99_143_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(203) is bound as output of CP function.
    -- CP-element group 204:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (4) 
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_update_start__ps
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_update_start_
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Update/req
      -- 
    req_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(204), ack => my_fetch4_99_143_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(204) is bound as output of CP function.
    -- CP-element group 205:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (4) 
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_sample_completed__ps
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Sample/ack
      -- 
    ack_814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch4_99_143_buf_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (4) 
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_update_completed__ps
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_my_fetch4_143_Update/ack
      -- 
    ack_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch4_99_143_buf_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (4) 
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_sample_start__ps
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Sample/req
      -- 
    req_831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(207), ack => n_fetch_val4_492_144_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(207) is bound as output of CP function.
    -- CP-element group 208:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (4) 
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_update_start__ps
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_update_start_
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Update/req
      -- 
    req_836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(208), ack => n_fetch_val4_492_144_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(208) is bound as output of CP function.
    -- CP-element group 209:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (4) 
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_sample_completed__ps
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Sample/ack
      -- 
    ack_832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val4_492_144_buf_ack_0, ack => access_T_CP_0_elements(209)); -- 
    -- CP-element group 210:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (4) 
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_update_completed__ps
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_fetch_val4_144_Update/ack
      -- 
    ack_837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val4_492_144_buf_ack_1, ack => access_T_CP_0_elements(210)); -- 
    -- CP-element group 211:  join  transition  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	30 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	33 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	32 
    -- CP-element group 211:  members (1) 
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_sample_start_
      -- 
    access_T_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33);
      gj_access_T_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  join  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	30 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	216 
    -- CP-element group 212: 	263 
    -- CP-element group 212: 	271 
    -- CP-element group 212: 	291 
    -- CP-element group 212: 	299 
    -- CP-element group 212: 	319 
    -- CP-element group 212: 	327 
    -- CP-element group 212: 	362 
    -- CP-element group 212: 	365 
    -- CP-element group 212: 	368 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	34 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_update_start_
      -- 
    access_T_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(216) & access_T_CP_0_elements(263) & access_T_CP_0_elements(271) & access_T_CP_0_elements(291) & access_T_CP_0_elements(299) & access_T_CP_0_elements(319) & access_T_CP_0_elements(327) & access_T_CP_0_elements(362) & access_T_CP_0_elements(365) & access_T_CP_0_elements(368);
      gj_access_T_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	32 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (1) 
      -- CP-element group 213: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_sample_start__ps
      -- 
    access_T_CP_0_elements(213) <= access_T_CP_0_elements(32);
    -- CP-element group 214:  join  transition  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	33 
    -- CP-element group 214:  members (1) 
      -- CP-element group 214: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(214) is bound as output of CP function.
    -- CP-element group 215:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	34 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_update_start__ps
      -- 
    access_T_CP_0_elements(215) <= access_T_CP_0_elements(34);
    -- CP-element group 216:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	35 
    -- CP-element group 216: 	31 
    -- CP-element group 216: 	261 
    -- CP-element group 216: 	269 
    -- CP-element group 216: 	289 
    -- CP-element group 216: 	297 
    -- CP-element group 216: 	317 
    -- CP-element group 216: 	325 
    -- CP-element group 216: 	361 
    -- CP-element group 216: 	364 
    -- CP-element group 216: 	367 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	212 
    -- CP-element group 216:  members (2) 
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(216) is bound as output of CP function.
    -- CP-element group 217:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	28 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_loopback_trigger
      -- 
    access_T_CP_0_elements(217) <= access_T_CP_0_elements(28);
    -- CP-element group 218:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_loopback_sample_req
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_loopback_sample_req_ps
      -- 
    phi_stmt_145_loopback_sample_req_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_145_loopback_sample_req_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(218), ack => phi_stmt_145_req_1); -- 
    -- Element group access_T_CP_0_elements(218) is bound as output of CP function.
    -- CP-element group 219:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	29 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_entry_trigger
      -- 
    access_T_CP_0_elements(219) <= access_T_CP_0_elements(29);
    -- CP-element group 220:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_entry_sample_req
      -- CP-element group 220: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_entry_sample_req_ps
      -- 
    phi_stmt_145_entry_sample_req_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_145_entry_sample_req_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(220), ack => phi_stmt_145_req_0); -- 
    -- Element group access_T_CP_0_elements(220) is bound as output of CP function.
    -- CP-element group 221:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (2) 
      -- CP-element group 221: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_phi_mux_ack
      -- CP-element group 221: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_145_phi_mux_ack_ps
      -- 
    phi_stmt_145_phi_mux_ack_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_145_ack_0, ack => access_T_CP_0_elements(221)); -- 
    -- CP-element group 222:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (4) 
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_sample_start__ps
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_sample_completed__ps
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(222) is bound as output of CP function.
    -- CP-element group 223:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_update_start__ps
      -- CP-element group 223: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_update_start_
      -- 
    -- Element group access_T_CP_0_elements(223) is bound as output of CP function.
    -- CP-element group 224:  join  transition  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	225 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (1) 
      -- CP-element group 224: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_update_completed__ps
      -- 
    access_T_CP_0_elements(224) <= access_T_CP_0_elements(225);
    -- CP-element group 225:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	224 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_148_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(225) is a control-delay.
    cp_element_225_delay: control_delay_element  generic map(name => " 225_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(223), ack => access_T_CP_0_elements(225), clk => clk, reset =>reset);
    -- CP-element group 226:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (4) 
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_sample_start__ps
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Sample/req
      -- 
    req_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(226), ack => n_row1_186_149_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(226) is bound as output of CP function.
    -- CP-element group 227:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (4) 
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_update_start__ps
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_update_start_
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Update/req
      -- 
    req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(227), ack => n_row1_186_149_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(227) is bound as output of CP function.
    -- CP-element group 228:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (4) 
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_sample_completed__ps
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Sample/ack
      -- 
    ack_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_186_149_buf_ack_0, ack => access_T_CP_0_elements(228)); -- 
    -- CP-element group 229:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (4) 
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_update_completed__ps
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row1_149_Update/ack
      -- 
    ack_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_186_149_buf_ack_1, ack => access_T_CP_0_elements(229)); -- 
    -- CP-element group 230:  join  transition  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	30 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	33 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	32 
    -- CP-element group 230:  members (1) 
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_sample_start_
      -- 
    access_T_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(33);
      gj_access_T_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	30 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	235 
    -- CP-element group 231: 	347 
    -- CP-element group 231: 	355 
    -- CP-element group 231: 	371 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	34 
    -- CP-element group 231:  members (1) 
      -- CP-element group 231: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_update_start_
      -- 
    access_T_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(235) & access_T_CP_0_elements(347) & access_T_CP_0_elements(355) & access_T_CP_0_elements(371);
      gj_access_T_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	32 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_sample_start__ps
      -- 
    access_T_CP_0_elements(232) <= access_T_CP_0_elements(32);
    -- CP-element group 233:  join  transition  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	33 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(233) is bound as output of CP function.
    -- CP-element group 234:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	34 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_update_start__ps
      -- 
    access_T_CP_0_elements(234) <= access_T_CP_0_elements(34);
    -- CP-element group 235:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	35 
    -- CP-element group 235: 	345 
    -- CP-element group 235: 	353 
    -- CP-element group 235: 	370 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	231 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(235) is bound as output of CP function.
    -- CP-element group 236:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	28 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_loopback_trigger
      -- 
    access_T_CP_0_elements(236) <= access_T_CP_0_elements(28);
    -- CP-element group 237:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_loopback_sample_req
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_loopback_sample_req_ps
      -- 
    phi_stmt_150_loopback_sample_req_892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_loopback_sample_req_892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(237), ack => phi_stmt_150_req_1); -- 
    -- Element group access_T_CP_0_elements(237) is bound as output of CP function.
    -- CP-element group 238:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	29 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (1) 
      -- CP-element group 238: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_entry_trigger
      -- 
    access_T_CP_0_elements(238) <= access_T_CP_0_elements(29);
    -- CP-element group 239:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_entry_sample_req
      -- CP-element group 239: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_entry_sample_req_ps
      -- 
    phi_stmt_150_entry_sample_req_895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_entry_sample_req_895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(239), ack => phi_stmt_150_req_0); -- 
    -- Element group access_T_CP_0_elements(239) is bound as output of CP function.
    -- CP-element group 240:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_phi_mux_ack
      -- CP-element group 240: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/phi_stmt_150_phi_mux_ack_ps
      -- 
    phi_stmt_150_phi_mux_ack_898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_150_ack_0, ack => access_T_CP_0_elements(240)); -- 
    -- CP-element group 241:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (4) 
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_sample_start__ps
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_sample_completed__ps
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(241) is bound as output of CP function.
    -- CP-element group 242:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_update_start__ps
      -- CP-element group 242: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_update_start_
      -- 
    -- Element group access_T_CP_0_elements(242) is bound as output of CP function.
    -- CP-element group 243:  join  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	244 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (1) 
      -- CP-element group 243: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_update_completed__ps
      -- 
    access_T_CP_0_elements(243) <= access_T_CP_0_elements(244);
    -- CP-element group 244:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	243 
    -- CP-element group 244:  members (1) 
      -- CP-element group 244: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_153_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(244) is a control-delay.
    cp_element_244_delay: control_delay_element  generic map(name => " 244_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(242), ack => access_T_CP_0_elements(244), clk => clk, reset =>reset);
    -- CP-element group 245:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (4) 
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_sample_start__ps
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Sample/req
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(245), ack => n_row2_194_154_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(245) is bound as output of CP function.
    -- CP-element group 246:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (4) 
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_update_start__ps
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_update_start_
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Update/req
      -- 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(246), ack => n_row2_194_154_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(246) is bound as output of CP function.
    -- CP-element group 247:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (4) 
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_sample_completed__ps
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Sample/ack
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_194_154_buf_ack_0, ack => access_T_CP_0_elements(247)); -- 
    -- CP-element group 248:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (4) 
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_update_completed__ps
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/R_n_row2_154_Update/ack
      -- 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_194_154_buf_ack_1, ack => access_T_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	30 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Sample/rr
      -- 
    rr_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(249), ack => type_cast_227_inst_req_0); -- 
    access_T_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(251);
      gj_access_T_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	33 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: 	257 
    -- CP-element group 250: 	263 
    -- CP-element group 250: 	271 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_update_start_
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Update/cr
      -- 
    cr_939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(250), ack => type_cast_227_inst_req_1); -- 
    access_T_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(252) & access_T_CP_0_elements(257) & access_T_CP_0_elements(263) & access_T_CP_0_elements(271);
      gj_access_T_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Sample/ra
      -- 
    ra_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_227_inst_ack_0, ack => access_T_CP_0_elements(251)); -- 
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	255 
    -- CP-element group 252: 	261 
    -- CP-element group 252: 	269 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	36 
    -- CP-element group 252: 	250 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_227_Update/ca
      -- 
    ca_940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_227_inst_ack_1, ack => access_T_CP_0_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	258 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	259 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	259 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_request/req
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_request/$entry
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_sample_start_
      -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(253), ack => addr_of_255_final_reg_req_0); -- 
    access_T_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(258) & access_T_CP_0_elements(259);
      gj_access_T_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	30 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	260 
    -- CP-element group 254: 	267 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	260 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_complete/$entry
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_complete/req
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_update_start_
      -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(254), ack => addr_of_255_final_reg_req_1); -- 
    access_T_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(260) & access_T_CP_0_elements(267);
      gj_access_T_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	121 
    -- CP-element group 255: 	41 
    -- CP-element group 255: 	252 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (13) 
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resized_1
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scaled_1
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_computed_1
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resize_1/$entry
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resize_1/$exit
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resize_1/index_resize_req
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_resize_1/index_resize_ack
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scale_1/$entry
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scale_1/$exit
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scale_1/scale_rename_req
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_index_scale_1/scale_rename_ack
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Sample/req
      -- 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(255), ack => array_obj_ref_254_index_offset_req_0); -- 
    access_T_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(121) & access_T_CP_0_elements(41) & access_T_CP_0_elements(252);
      gj_access_T_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	30 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: 	259 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_update_start
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Update/req
      -- 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(256), ack => array_obj_ref_254_index_offset_req_1); -- 
    access_T_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(258) & access_T_CP_0_elements(259);
      gj_access_T_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	374 
    -- CP-element group 257: marked-successors 
    -- CP-element group 257: 	117 
    -- CP-element group 257: 	37 
    -- CP-element group 257: 	250 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_sample_complete
      -- CP-element group 257: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Sample/ack
      -- 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_254_index_offset_ack_0, ack => access_T_CP_0_elements(257)); -- 
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	253 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (8) 
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_base_plus_offset/sum_rename_ack
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_base_plus_offset/sum_rename_req
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_base_plus_offset/$exit
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_base_plus_offset/$entry
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_root_address_calculated
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_offset_calculated
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_254_final_index_sum_regn_Update/ack
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_254_index_offset_ack_1, ack => access_T_CP_0_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	253 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	253 
    -- CP-element group 259: 	256 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_request/ack
      -- CP-element group 259: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_request/$exit
      -- CP-element group 259: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_sample_completed_
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_255_final_reg_ack_0, ack => access_T_CP_0_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	254 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	265 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	254 
    -- CP-element group 260:  members (19) 
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_complete/$exit
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_addrgen/root_register_ack
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_addrgen/root_register_req
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_addrgen/$exit
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_addrgen/$entry
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_plus_offset/sum_rename_ack
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_complete/ack
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_plus_offset/sum_rename_req
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_plus_offset/$exit
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_plus_offset/$entry
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_addr_resize/base_resize_ack
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_addr_resize/base_resize_req
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_addr_resize/$exit
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_addr_resize/$entry
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_address_resized
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_root_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_word_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_base_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_255_update_completed_
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_255_final_reg_ack_1, ack => access_T_CP_0_elements(260)); -- 
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	121 
    -- CP-element group 261: 	41 
    -- CP-element group 261: 	216 
    -- CP-element group 261: 	252 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Sample/req
      -- CP-element group 261: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Sample/$entry
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(261), ack => W_fn1_254_delayed_7_0_257_inst_req_0); -- 
    access_T_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(121) & access_T_CP_0_elements(41) & access_T_CP_0_elements(216) & access_T_CP_0_elements(252) & access_T_CP_0_elements(263);
      gj_access_T_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	264 
    -- CP-element group 262: 	267 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_update_start_
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Update/req
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Update/$entry
      -- 
    req_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(262), ack => W_fn1_254_delayed_7_0_257_inst_req_1); -- 
    access_T_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(264) & access_T_CP_0_elements(267);
      gj_access_T_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	117 
    -- CP-element group 263: 	37 
    -- CP-element group 263: 	212 
    -- CP-element group 263: 	250 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Sample/$exit
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_254_delayed_7_0_257_inst_ack_0, ack => access_T_CP_0_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_259_update_completed_
      -- 
    ack_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_254_delayed_7_0_257_inst_ack_1, ack => access_T_CP_0_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	260 
    -- CP-element group 265: 	264 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (5) 
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/word_0/rr
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/word_0/$entry
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/$entry
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_sample_start_
      -- 
    rr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(265), ack => ptr_deref_263_load_0_req_0); -- 
    access_T_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(260) & access_T_CP_0_elements(264) & access_T_CP_0_elements(267);
      gj_access_T_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	33 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (5) 
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/word_0/cr
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/word_0/$entry
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/$entry
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_update_start_
      -- 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(266), ack => ptr_deref_263_load_0_req_1); -- 
    access_T_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(268);
      gj_access_T_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	254 
    -- CP-element group 267: 	262 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (5) 
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/word_0/ra
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/word_0/$exit
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/word_access_start/$exit
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_sample_completed_
      -- 
    ra_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_load_0_ack_0, ack => access_T_CP_0_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	374 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	135 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (9) 
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/ptr_deref_263_Merge/merge_req
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/ptr_deref_263_Merge/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/ptr_deref_263_Merge/$entry
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/word_0/ca
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/word_0/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/word_access_complete/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_263_Update/ptr_deref_263_Merge/merge_ack
      -- 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_load_0_ack_1, ack => access_T_CP_0_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	121 
    -- CP-element group 269: 	41 
    -- CP-element group 269: 	216 
    -- CP-element group 269: 	252 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Sample/req
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_sample_start_
      -- 
    req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(269), ack => W_fn1_260_delayed_13_0_265_inst_req_0); -- 
    access_T_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(121) & access_T_CP_0_elements(41) & access_T_CP_0_elements(216) & access_T_CP_0_elements(252) & access_T_CP_0_elements(271);
      gj_access_T_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	33 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Update/req
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_update_start_
      -- 
    req_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(270), ack => W_fn1_260_delayed_13_0_265_inst_req_1); -- 
    access_T_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(272);
      gj_access_T_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	117 
    -- CP-element group 271: 	37 
    -- CP-element group 271: 	212 
    -- CP-element group 271: 	250 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_sample_completed_
      -- 
    ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_260_delayed_13_0_265_inst_ack_0, ack => access_T_CP_0_elements(271)); -- 
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	374 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	135 
    -- CP-element group 272: 	270 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_267_update_completed_
      -- 
    ack_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_260_delayed_13_0_265_inst_ack_1, ack => access_T_CP_0_elements(272)); -- 
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	140 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Sample/req
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_sample_start_
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(273), ack => W_fetch_val1_262_delayed_13_0_268_inst_req_0); -- 
    access_T_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(140) & access_T_CP_0_elements(275);
      gj_access_T_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	33 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Update/req
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_update_start_
      -- 
    req_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(274), ack => W_fetch_val1_262_delayed_13_0_268_inst_req_1); -- 
    access_T_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(276);
      gj_access_T_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	136 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_sample_completed_
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val1_262_delayed_13_0_268_inst_ack_0, ack => access_T_CP_0_elements(275)); -- 
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	374 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	135 
    -- CP-element group 276: 	274 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_270_update_completed_
      -- 
    ack_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val1_262_delayed_13_0_268_inst_ack_1, ack => access_T_CP_0_elements(276)); -- 
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	30 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_sample_start_
      -- CP-element group 277: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Sample/rr
      -- CP-element group 277: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Sample/$entry
      -- 
    rr_1086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(277), ack => type_cast_299_inst_req_0); -- 
    access_T_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(279);
      gj_access_T_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	33 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: 	285 
    -- CP-element group 278: 	291 
    -- CP-element group 278: 	299 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Update/cr
      -- CP-element group 278: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Update/$entry
      -- CP-element group 278: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_update_start_
      -- 
    cr_1091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(278), ack => type_cast_299_inst_req_1); -- 
    access_T_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(280) & access_T_CP_0_elements(285) & access_T_CP_0_elements(291) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_sample_completed_
      -- 
    ra_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_299_inst_ack_0, ack => access_T_CP_0_elements(279)); -- 
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280: 	289 
    -- CP-element group 280: 	297 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	55 
    -- CP-element group 280: 	278 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Update/ca
      -- CP-element group 280: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_299_update_completed_
      -- 
    ca_1092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_299_inst_ack_1, ack => access_T_CP_0_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	286 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	287 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	287 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_request/req
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_request/$entry
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_sample_start_
      -- 
    req_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(281), ack => addr_of_327_final_reg_req_0); -- 
    access_T_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(286) & access_T_CP_0_elements(287);
      gj_access_T_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	30 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	288 
    -- CP-element group 282: 	295 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	288 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_complete/req
      -- CP-element group 282: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_complete/$entry
      -- CP-element group 282: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_update_start_
      -- 
    req_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(282), ack => addr_of_327_final_reg_req_1); -- 
    access_T_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(288) & access_T_CP_0_elements(295);
      gj_access_T_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	121 
    -- CP-element group 283: 	60 
    -- CP-element group 283: 	280 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (13) 
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resized_1
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scale_1/scale_rename_ack
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scale_1/scale_rename_req
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scale_1/$exit
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scale_1/$entry
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resize_1/index_resize_ack
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resize_1/index_resize_req
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resize_1/$exit
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_resize_1/$entry
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_computed_1
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_index_scaled_1
      -- 
    req_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(283), ack => array_obj_ref_326_index_offset_req_0); -- 
    access_T_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(121) & access_T_CP_0_elements(60) & access_T_CP_0_elements(280);
      gj_access_T_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	30 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	286 
    -- CP-element group 284: 	287 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_update_start
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Update/req
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Update/$entry
      -- 
    req_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(284), ack => array_obj_ref_326_index_offset_req_1); -- 
    access_T_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(286) & access_T_CP_0_elements(287);
      gj_access_T_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	374 
    -- CP-element group 285: marked-successors 
    -- CP-element group 285: 	117 
    -- CP-element group 285: 	56 
    -- CP-element group 285: 	278 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_sample_complete
      -- 
    ack_1118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_326_index_offset_ack_0, ack => access_T_CP_0_elements(285)); -- 
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	281 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	284 
    -- CP-element group 286:  members (8) 
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_offset_calculated
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_root_address_calculated
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_base_plus_offset/sum_rename_ack
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_base_plus_offset/sum_rename_req
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_base_plus_offset/$exit
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_base_plus_offset/$entry
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_326_final_index_sum_regn_Update/$exit
      -- 
    ack_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_326_index_offset_ack_1, ack => access_T_CP_0_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	281 
    -- CP-element group 287: successors 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	281 
    -- CP-element group 287: 	284 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_request/ack
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_request/$exit
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_sample_completed_
      -- 
    ack_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_327_final_reg_ack_0, ack => access_T_CP_0_elements(287)); -- 
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	282 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	293 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	282 
    -- CP-element group 288:  members (19) 
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_complete/ack
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_complete/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_addrgen/root_register_ack
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_addrgen/root_register_req
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_327_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_plus_offset/sum_rename_req
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_addrgen/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_addrgen/$entry
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_plus_offset/sum_rename_ack
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_plus_offset/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_plus_offset/$entry
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_addr_resize/base_resize_ack
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_addr_resize/base_resize_req
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_addr_resize/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_addr_resize/$entry
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_address_resized
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_root_address_calculated
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_word_address_calculated
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_base_address_calculated
      -- 
    ack_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_327_final_reg_ack_1, ack => access_T_CP_0_elements(288)); -- 
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	121 
    -- CP-element group 289: 	60 
    -- CP-element group 289: 	216 
    -- CP-element group 289: 	280 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Sample/req
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_sample_start_
      -- 
    req_1146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(289), ack => W_fn2_314_delayed_7_0_329_inst_req_0); -- 
    access_T_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(121) & access_T_CP_0_elements(60) & access_T_CP_0_elements(216) & access_T_CP_0_elements(280) & access_T_CP_0_elements(291);
      gj_access_T_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: 	295 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_update_start_
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Update/req
      -- 
    req_1151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(290), ack => W_fn2_314_delayed_7_0_329_inst_req_1); -- 
    access_T_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(292) & access_T_CP_0_elements(295);
      gj_access_T_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	117 
    -- CP-element group 291: 	56 
    -- CP-element group 291: 	212 
    -- CP-element group 291: 	278 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_sample_completed_
      -- 
    ack_1147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_314_delayed_7_0_329_inst_ack_0, ack => access_T_CP_0_elements(291)); -- 
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	290 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_331_Update/ack
      -- 
    ack_1152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_314_delayed_7_0_329_inst_ack_1, ack => access_T_CP_0_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	288 
    -- CP-element group 293: 	292 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (5) 
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/word_0/rr
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/word_0/$entry
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/$entry
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/$entry
      -- 
    rr_1185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(293), ack => ptr_deref_335_load_0_req_0); -- 
    access_T_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(288) & access_T_CP_0_elements(292) & access_T_CP_0_elements(295);
      gj_access_T_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	33 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (5) 
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_update_start_
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/word_0/cr
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/word_0/$entry
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/$entry
      -- 
    cr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(294), ack => ptr_deref_335_load_0_req_1); -- 
    access_T_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(296);
      gj_access_T_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	282 
    -- CP-element group 295: 	290 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (5) 
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/word_0/ra
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/word_0/$exit
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/word_access_start/$exit
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Sample/$exit
      -- 
    ra_1186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_335_load_0_ack_0, ack => access_T_CP_0_elements(295)); -- 
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	374 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	154 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (9) 
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/word_0/ca
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/word_0/$exit
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/word_access_complete/$exit
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/ptr_deref_335_Merge/merge_ack
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/ptr_deref_335_Merge/merge_req
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/ptr_deref_335_Merge/$exit
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_Update/ptr_deref_335_Merge/$entry
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_335_update_completed_
      -- 
    ca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_335_load_0_ack_1, ack => access_T_CP_0_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	121 
    -- CP-element group 297: 	60 
    -- CP-element group 297: 	216 
    -- CP-element group 297: 	280 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Sample/req
      -- CP-element group 297: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_sample_start_
      -- 
    req_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(297), ack => W_fn2_320_delayed_13_0_337_inst_req_0); -- 
    access_T_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(121) & access_T_CP_0_elements(60) & access_T_CP_0_elements(216) & access_T_CP_0_elements(280) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	33 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Update/req
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_update_start_
      -- 
    req_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(298), ack => W_fn2_320_delayed_13_0_337_inst_req_1); -- 
    access_T_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(300);
      gj_access_T_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	117 
    -- CP-element group 299: 	56 
    -- CP-element group 299: 	212 
    -- CP-element group 299: 	278 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_sample_completed_
      -- 
    ack_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_320_delayed_13_0_337_inst_ack_0, ack => access_T_CP_0_elements(299)); -- 
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	374 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	154 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_339_Update/ack
      -- 
    ack_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_320_delayed_13_0_337_inst_ack_1, ack => access_T_CP_0_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	159 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Sample/req
      -- CP-element group 301: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_sample_start_
      -- 
    req_1224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(301), ack => W_fetch_val2_322_delayed_13_0_340_inst_req_0); -- 
    access_T_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(159) & access_T_CP_0_elements(303);
      gj_access_T_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	33 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Update/req
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_update_start_
      -- 
    req_1229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(302), ack => W_fetch_val2_322_delayed_13_0_340_inst_req_1); -- 
    access_T_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(304);
      gj_access_T_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	155 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_sample_completed_
      -- 
    ack_1225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val2_322_delayed_13_0_340_inst_ack_0, ack => access_T_CP_0_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	374 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	154 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_342_update_completed_
      -- 
    ack_1230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val2_322_delayed_13_0_340_inst_ack_1, ack => access_T_CP_0_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	30 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Sample/rr
      -- 
    rr_1238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(305), ack => type_cast_371_inst_req_0); -- 
    access_T_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(307);
      gj_access_T_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	33 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: 	313 
    -- CP-element group 306: 	319 
    -- CP-element group 306: 	327 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_update_start_
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Update/cr
      -- 
    cr_1243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(306), ack => type_cast_371_inst_req_1); -- 
    access_T_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(308) & access_T_CP_0_elements(313) & access_T_CP_0_elements(319) & access_T_CP_0_elements(327);
      gj_access_T_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Sample/ra
      -- 
    ra_1239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_0, ack => access_T_CP_0_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	311 
    -- CP-element group 308: 	317 
    -- CP-element group 308: 	325 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	76 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_371_Update/ca
      -- 
    ca_1244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_371_inst_ack_1, ack => access_T_CP_0_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	314 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	315 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	315 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_request/$entry
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_request/req
      -- 
    req_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(309), ack => addr_of_399_final_reg_req_0); -- 
    access_T_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(314) & access_T_CP_0_elements(315);
      gj_access_T_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	30 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	316 
    -- CP-element group 310: 	323 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	316 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_update_start_
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_complete/$entry
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_complete/req
      -- 
    req_1289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(310), ack => addr_of_399_final_reg_req_1); -- 
    access_T_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(316) & access_T_CP_0_elements(323);
      gj_access_T_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	79 
    -- CP-element group 311: 	121 
    -- CP-element group 311: 	308 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311:  members (13) 
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resized_1
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scaled_1
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_computed_1
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resize_1/$entry
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resize_1/$exit
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resize_1/index_resize_req
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_resize_1/index_resize_ack
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scale_1/$entry
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scale_1/$exit
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scale_1/scale_rename_req
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_index_scale_1/scale_rename_ack
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Sample/req
      -- 
    req_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(311), ack => array_obj_ref_398_index_offset_req_0); -- 
    access_T_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(79) & access_T_CP_0_elements(121) & access_T_CP_0_elements(308);
      gj_access_T_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	30 
    -- CP-element group 312: marked-predecessors 
    -- CP-element group 312: 	314 
    -- CP-element group 312: 	315 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	314 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_update_start
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Update/req
      -- 
    req_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(312), ack => array_obj_ref_398_index_offset_req_1); -- 
    access_T_cp_element_group_312: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_312"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(314) & access_T_CP_0_elements(315);
      gj_access_T_cp_element_group_312 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(312), clk => clk, reset => reset); --
    end block;
    -- CP-element group 313:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	311 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	374 
    -- CP-element group 313: marked-successors 
    -- CP-element group 313: 	77 
    -- CP-element group 313: 	117 
    -- CP-element group 313: 	306 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_sample_complete
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Sample/ack
      -- 
    ack_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_398_index_offset_ack_0, ack => access_T_CP_0_elements(313)); -- 
    -- CP-element group 314:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	312 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	309 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	312 
    -- CP-element group 314:  members (8) 
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_root_address_calculated
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_offset_calculated
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_final_index_sum_regn_Update/ack
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_base_plus_offset/$entry
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_base_plus_offset/$exit
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_base_plus_offset/sum_rename_req
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_398_base_plus_offset/sum_rename_ack
      -- 
    ack_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_398_index_offset_ack_1, ack => access_T_CP_0_elements(314)); -- 
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	309 
    -- CP-element group 315: successors 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	309 
    -- CP-element group 315: 	312 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_request/$exit
      -- CP-element group 315: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_request/ack
      -- 
    ack_1285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_399_final_reg_ack_0, ack => access_T_CP_0_elements(315)); -- 
    -- CP-element group 316:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	310 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	321 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	310 
    -- CP-element group 316:  members (19) 
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_complete/$exit
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_399_complete/ack
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_root_address_calculated
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_address_resized
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_addr_resize/$entry
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_addr_resize/$exit
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_addr_resize/base_resize_req
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_addr_resize/base_resize_ack
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_plus_offset/$entry
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_plus_offset/$exit
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_plus_offset/sum_rename_req
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_base_plus_offset/sum_rename_ack
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_addrgen/$entry
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_addrgen/$exit
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_addrgen/root_register_req
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_word_addrgen/root_register_ack
      -- 
    ack_1290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_399_final_reg_ack_1, ack => access_T_CP_0_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	79 
    -- CP-element group 317: 	121 
    -- CP-element group 317: 	216 
    -- CP-element group 317: 	308 
    -- CP-element group 317: marked-predecessors 
    -- CP-element group 317: 	319 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Sample/req
      -- 
    req_1298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(317), ack => W_fn3_374_delayed_7_0_401_inst_req_0); -- 
    access_T_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(79) & access_T_CP_0_elements(121) & access_T_CP_0_elements(216) & access_T_CP_0_elements(308) & access_T_CP_0_elements(319);
      gj_access_T_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	320 
    -- CP-element group 318: 	323 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_update_start_
      -- CP-element group 318: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Update/req
      -- 
    req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(318), ack => W_fn3_374_delayed_7_0_401_inst_req_1); -- 
    access_T_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(320) & access_T_CP_0_elements(323);
      gj_access_T_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: successors 
    -- CP-element group 319: marked-successors 
    -- CP-element group 319: 	77 
    -- CP-element group 319: 	117 
    -- CP-element group 319: 	212 
    -- CP-element group 319: 	306 
    -- CP-element group 319: 	317 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Sample/ack
      -- 
    ack_1299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_374_delayed_7_0_401_inst_ack_0, ack => access_T_CP_0_elements(319)); -- 
    -- CP-element group 320:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	318 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_403_Update/ack
      -- 
    ack_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_374_delayed_7_0_401_inst_ack_1, ack => access_T_CP_0_elements(320)); -- 
    -- CP-element group 321:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	316 
    -- CP-element group 321: 	320 
    -- CP-element group 321: marked-predecessors 
    -- CP-element group 321: 	323 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (5) 
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_sample_start_
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/$entry
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/$entry
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/word_0/$entry
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/word_0/rr
      -- 
    rr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(321), ack => ptr_deref_407_load_0_req_0); -- 
    access_T_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(316) & access_T_CP_0_elements(320) & access_T_CP_0_elements(323);
      gj_access_T_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	33 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (5) 
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_update_start_
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/$entry
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/$entry
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/word_0/$entry
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/word_0/cr
      -- 
    cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(322), ack => ptr_deref_407_load_0_req_1); -- 
    access_T_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(324);
      gj_access_T_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: successors 
    -- CP-element group 323: marked-successors 
    -- CP-element group 323: 	310 
    -- CP-element group 323: 	318 
    -- CP-element group 323: 	321 
    -- CP-element group 323:  members (5) 
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/$exit
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/word_0/$exit
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Sample/word_access_start/word_0/ra
      -- 
    ra_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_407_load_0_ack_0, ack => access_T_CP_0_elements(323)); -- 
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	374 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	173 
    -- CP-element group 324: 	322 
    -- CP-element group 324:  members (9) 
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/$exit
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/word_0/$exit
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/word_access_complete/word_0/ca
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/ptr_deref_407_Merge/$entry
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/ptr_deref_407_Merge/$exit
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/ptr_deref_407_Merge/merge_req
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_407_Update/ptr_deref_407_Merge/merge_ack
      -- 
    ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_407_load_0_ack_1, ack => access_T_CP_0_elements(324)); -- 
    -- CP-element group 325:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	79 
    -- CP-element group 325: 	121 
    -- CP-element group 325: 	216 
    -- CP-element group 325: 	308 
    -- CP-element group 325: marked-predecessors 
    -- CP-element group 325: 	327 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Sample/req
      -- 
    req_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(325), ack => W_fn3_380_delayed_13_0_409_inst_req_0); -- 
    access_T_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(79) & access_T_CP_0_elements(121) & access_T_CP_0_elements(216) & access_T_CP_0_elements(308) & access_T_CP_0_elements(327);
      gj_access_T_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	33 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_update_start_
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Update/req
      -- 
    req_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(326), ack => W_fn3_380_delayed_13_0_409_inst_req_1); -- 
    access_T_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(328);
      gj_access_T_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: marked-successors 
    -- CP-element group 327: 	77 
    -- CP-element group 327: 	117 
    -- CP-element group 327: 	212 
    -- CP-element group 327: 	306 
    -- CP-element group 327: 	325 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Sample/ack
      -- 
    ack_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_380_delayed_13_0_409_inst_ack_0, ack => access_T_CP_0_elements(327)); -- 
    -- CP-element group 328:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	374 
    -- CP-element group 328: marked-successors 
    -- CP-element group 328: 	173 
    -- CP-element group 328: 	326 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_411_Update/ack
      -- 
    ack_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_380_delayed_13_0_409_inst_ack_1, ack => access_T_CP_0_elements(328)); -- 
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	178 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_sample_start_
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Sample/req
      -- 
    req_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(329), ack => W_fetch_val3_382_delayed_13_0_412_inst_req_0); -- 
    access_T_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(178) & access_T_CP_0_elements(331);
      gj_access_T_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	33 
    -- CP-element group 330: marked-predecessors 
    -- CP-element group 330: 	332 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_update_start_
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Update/req
      -- 
    req_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(330), ack => W_fetch_val3_382_delayed_13_0_412_inst_req_1); -- 
    access_T_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(332);
      gj_access_T_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	174 
    -- CP-element group 331: 	329 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Sample/ack
      -- 
    ack_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val3_382_delayed_13_0_412_inst_ack_0, ack => access_T_CP_0_elements(331)); -- 
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	374 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	173 
    -- CP-element group 332: 	330 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_414_Update/ack
      -- 
    ack_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val3_382_delayed_13_0_412_inst_ack_1, ack => access_T_CP_0_elements(332)); -- 
    -- CP-element group 333:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	30 
    -- CP-element group 333: marked-predecessors 
    -- CP-element group 333: 	335 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Sample/rr
      -- 
    rr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(333), ack => type_cast_443_inst_req_0); -- 
    access_T_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(335);
      gj_access_T_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	33 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: 	341 
    -- CP-element group 334: 	347 
    -- CP-element group 334: 	355 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_update_start_
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Update/cr
      -- 
    cr_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(334), ack => type_cast_443_inst_req_1); -- 
    access_T_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(336) & access_T_CP_0_elements(341) & access_T_CP_0_elements(347) & access_T_CP_0_elements(355);
      gj_access_T_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: successors 
    -- CP-element group 335: marked-successors 
    -- CP-element group 335: 	333 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Sample/ra
      -- 
    ra_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_0, ack => access_T_CP_0_elements(335)); -- 
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	339 
    -- CP-element group 336: 	345 
    -- CP-element group 336: 	353 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	95 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/type_cast_443_Update/ca
      -- 
    ca_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_443_inst_ack_1, ack => access_T_CP_0_elements(336)); -- 
    -- CP-element group 337:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	342 
    -- CP-element group 337: marked-predecessors 
    -- CP-element group 337: 	343 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	343 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_request/$entry
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_request/req
      -- 
    req_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(337), ack => addr_of_471_final_reg_req_0); -- 
    access_T_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(342) & access_T_CP_0_elements(343);
      gj_access_T_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	30 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	344 
    -- CP-element group 338: 	351 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	344 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_update_start_
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_complete/$entry
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_complete/req
      -- 
    req_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(338), ack => addr_of_471_final_reg_req_1); -- 
    access_T_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(344) & access_T_CP_0_elements(351);
      gj_access_T_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	100 
    -- CP-element group 339: 	121 
    -- CP-element group 339: 	336 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (13) 
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resized_1
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scaled_1
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_computed_1
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resize_1/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resize_1/$exit
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resize_1/index_resize_req
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_resize_1/index_resize_ack
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scale_1/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scale_1/$exit
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scale_1/scale_rename_req
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_index_scale_1/scale_rename_ack
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Sample/req
      -- 
    req_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(339), ack => array_obj_ref_470_index_offset_req_0); -- 
    access_T_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(100) & access_T_CP_0_elements(121) & access_T_CP_0_elements(336);
      gj_access_T_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	30 
    -- CP-element group 340: marked-predecessors 
    -- CP-element group 340: 	342 
    -- CP-element group 340: 	343 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	342 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_update_start
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Update/$entry
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Update/req
      -- 
    req_1426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(340), ack => array_obj_ref_470_index_offset_req_1); -- 
    access_T_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(30) & access_T_CP_0_elements(342) & access_T_CP_0_elements(343);
      gj_access_T_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	374 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	96 
    -- CP-element group 341: 	117 
    -- CP-element group 341: 	334 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_sample_complete
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Sample/ack
      -- 
    ack_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_470_index_offset_ack_0, ack => access_T_CP_0_elements(341)); -- 
    -- CP-element group 342:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	337 
    -- CP-element group 342: marked-successors 
    -- CP-element group 342: 	340 
    -- CP-element group 342:  members (8) 
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_root_address_calculated
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_offset_calculated
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_final_index_sum_regn_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_base_plus_offset/$entry
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_base_plus_offset/$exit
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_base_plus_offset/sum_rename_req
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/array_obj_ref_470_base_plus_offset/sum_rename_ack
      -- 
    ack_1427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_470_index_offset_ack_1, ack => access_T_CP_0_elements(342)); -- 
    -- CP-element group 343:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	337 
    -- CP-element group 343: successors 
    -- CP-element group 343: marked-successors 
    -- CP-element group 343: 	337 
    -- CP-element group 343: 	340 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_request/$exit
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_request/ack
      -- 
    ack_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_471_final_reg_ack_0, ack => access_T_CP_0_elements(343)); -- 
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	338 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	349 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	338 
    -- CP-element group 344:  members (19) 
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_complete/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/addr_of_471_complete/ack
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_address_calculated
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_address_calculated
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_root_address_calculated
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_address_resized
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_addr_resize/$entry
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_addr_resize/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_addr_resize/base_resize_req
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_addr_resize/base_resize_ack
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_plus_offset/$entry
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_plus_offset/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_plus_offset/sum_rename_req
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_base_plus_offset/sum_rename_ack
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_addrgen/$entry
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_addrgen/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_addrgen/root_register_req
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_word_addrgen/root_register_ack
      -- 
    ack_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_471_final_reg_ack_1, ack => access_T_CP_0_elements(344)); -- 
    -- CP-element group 345:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	100 
    -- CP-element group 345: 	121 
    -- CP-element group 345: 	235 
    -- CP-element group 345: 	336 
    -- CP-element group 345: marked-predecessors 
    -- CP-element group 345: 	347 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_sample_start_
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Sample/req
      -- 
    req_1450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(345), ack => W_fn4_434_delayed_7_0_473_inst_req_0); -- 
    access_T_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(100) & access_T_CP_0_elements(121) & access_T_CP_0_elements(235) & access_T_CP_0_elements(336) & access_T_CP_0_elements(347);
      gj_access_T_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: 	351 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_update_start_
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Update/req
      -- 
    req_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(346), ack => W_fn4_434_delayed_7_0_473_inst_req_1); -- 
    access_T_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(348) & access_T_CP_0_elements(351);
      gj_access_T_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: marked-successors 
    -- CP-element group 347: 	96 
    -- CP-element group 347: 	117 
    -- CP-element group 347: 	231 
    -- CP-element group 347: 	334 
    -- CP-element group 347: 	345 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Sample/ack
      -- 
    ack_1451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn4_434_delayed_7_0_473_inst_ack_0, ack => access_T_CP_0_elements(347)); -- 
    -- CP-element group 348:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348: marked-successors 
    -- CP-element group 348: 	346 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_475_Update/ack
      -- 
    ack_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn4_434_delayed_7_0_473_inst_ack_1, ack => access_T_CP_0_elements(348)); -- 
    -- CP-element group 349:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	344 
    -- CP-element group 349: 	348 
    -- CP-element group 349: marked-predecessors 
    -- CP-element group 349: 	351 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (5) 
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/$entry
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/word_0/$entry
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/word_0/rr
      -- 
    rr_1489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(349), ack => ptr_deref_479_load_0_req_0); -- 
    access_T_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(344) & access_T_CP_0_elements(348) & access_T_CP_0_elements(351);
      gj_access_T_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	33 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	352 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (5) 
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_update_start_
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/word_0/$entry
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/word_0/cr
      -- 
    cr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(350), ack => ptr_deref_479_load_0_req_1); -- 
    access_T_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(352);
      gj_access_T_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: successors 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	338 
    -- CP-element group 351: 	346 
    -- CP-element group 351: 	349 
    -- CP-element group 351:  members (5) 
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_sample_completed_
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/$exit
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/word_0/$exit
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Sample/word_access_start/word_0/ra
      -- 
    ra_1490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_479_load_0_ack_0, ack => access_T_CP_0_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	374 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	192 
    -- CP-element group 352: 	350 
    -- CP-element group 352:  members (9) 
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_update_completed_
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/word_0/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/word_access_complete/word_0/ca
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/ptr_deref_479_Merge/$entry
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/ptr_deref_479_Merge/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/ptr_deref_479_Merge/merge_req
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/ptr_deref_479_Update/ptr_deref_479_Merge/merge_ack
      -- 
    ca_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_479_load_0_ack_1, ack => access_T_CP_0_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	100 
    -- CP-element group 353: 	121 
    -- CP-element group 353: 	235 
    -- CP-element group 353: 	336 
    -- CP-element group 353: marked-predecessors 
    -- CP-element group 353: 	355 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Sample/req
      -- 
    req_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(353), ack => W_fn4_440_delayed_13_0_481_inst_req_0); -- 
    access_T_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(100) & access_T_CP_0_elements(121) & access_T_CP_0_elements(235) & access_T_CP_0_elements(336) & access_T_CP_0_elements(355);
      gj_access_T_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	33 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_update_start_
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Update/$entry
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Update/req
      -- 
    req_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(354), ack => W_fn4_440_delayed_13_0_481_inst_req_1); -- 
    access_T_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(356);
      gj_access_T_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: marked-successors 
    -- CP-element group 355: 	96 
    -- CP-element group 355: 	117 
    -- CP-element group 355: 	231 
    -- CP-element group 355: 	334 
    -- CP-element group 355: 	353 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Sample/ack
      -- 
    ack_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn4_440_delayed_13_0_481_inst_ack_0, ack => access_T_CP_0_elements(355)); -- 
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	374 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	192 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_483_Update/ack
      -- 
    ack_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn4_440_delayed_13_0_481_inst_ack_1, ack => access_T_CP_0_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	197 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	359 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Sample/req
      -- 
    req_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(357), ack => W_fetch_val4_442_delayed_13_0_484_inst_req_0); -- 
    access_T_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(197) & access_T_CP_0_elements(359);
      gj_access_T_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	33 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_update_start_
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Update/$entry
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Update/req
      -- 
    req_1533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(358), ack => W_fetch_val4_442_delayed_13_0_484_inst_req_1); -- 
    access_T_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(360);
      gj_access_T_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: marked-successors 
    -- CP-element group 359: 	193 
    -- CP-element group 359: 	357 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Sample/ack
      -- 
    ack_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val4_442_delayed_13_0_484_inst_ack_0, ack => access_T_CP_0_elements(359)); -- 
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	374 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	192 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/assign_stmt_486_Update/ack
      -- 
    ack_1534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val4_442_delayed_13_0_484_inst_ack_1, ack => access_T_CP_0_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	41 
    -- CP-element group 361: 	140 
    -- CP-element group 361: 	216 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	363 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_sample_start_
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Sample/req
      -- 
    req_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(361), ack => WPIPE_input_pipe1_494_inst_req_0); -- 
    access_T_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(41) & access_T_CP_0_elements(140) & access_T_CP_0_elements(216) & access_T_CP_0_elements(363);
      gj_access_T_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362: marked-successors 
    -- CP-element group 362: 	136 
    -- CP-element group 362: 	37 
    -- CP-element group 362: 	212 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_sample_completed_
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_update_start_
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Sample/ack
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Update/$entry
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Update/req
      -- 
    ack_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_494_inst_ack_0, ack => access_T_CP_0_elements(362)); -- 
    req_1547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(362), ack => WPIPE_input_pipe1_494_inst_req_1); -- 
    -- CP-element group 363:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	374 
    -- CP-element group 363: marked-successors 
    -- CP-element group 363: 	361 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_update_completed_
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe1_494_Update/ack
      -- 
    ack_1548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_494_inst_ack_1, ack => access_T_CP_0_elements(363)); -- 
    -- CP-element group 364:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	60 
    -- CP-element group 364: 	159 
    -- CP-element group 364: 	216 
    -- CP-element group 364: marked-predecessors 
    -- CP-element group 364: 	366 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_sample_start_
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Sample/$entry
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Sample/req
      -- 
    req_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(364), ack => WPIPE_input_pipe2_498_inst_req_0); -- 
    access_T_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(60) & access_T_CP_0_elements(159) & access_T_CP_0_elements(216) & access_T_CP_0_elements(366);
      gj_access_T_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	56 
    -- CP-element group 365: 	155 
    -- CP-element group 365: 	212 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_update_start_
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Sample/ack
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Update/req
      -- 
    ack_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_498_inst_ack_0, ack => access_T_CP_0_elements(365)); -- 
    req_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(365), ack => WPIPE_input_pipe2_498_inst_req_1); -- 
    -- CP-element group 366:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	374 
    -- CP-element group 366: marked-successors 
    -- CP-element group 366: 	364 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe2_498_Update/ack
      -- 
    ack_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_498_inst_ack_1, ack => access_T_CP_0_elements(366)); -- 
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	79 
    -- CP-element group 367: 	178 
    -- CP-element group 367: 	216 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_sample_start_
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Sample/req
      -- 
    req_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(367), ack => WPIPE_input_pipe3_502_inst_req_0); -- 
    access_T_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(79) & access_T_CP_0_elements(178) & access_T_CP_0_elements(216) & access_T_CP_0_elements(369);
      gj_access_T_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	77 
    -- CP-element group 368: 	174 
    -- CP-element group 368: 	212 
    -- CP-element group 368:  members (6) 
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_update_start_
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Sample/ack
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Update/req
      -- 
    ack_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_502_inst_ack_0, ack => access_T_CP_0_elements(368)); -- 
    req_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(368), ack => WPIPE_input_pipe3_502_inst_req_1); -- 
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe3_502_Update/ack
      -- 
    ack_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_502_inst_ack_1, ack => access_T_CP_0_elements(369)); -- 
    -- CP-element group 370:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	100 
    -- CP-element group 370: 	197 
    -- CP-element group 370: 	235 
    -- CP-element group 370: marked-predecessors 
    -- CP-element group 370: 	372 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Sample/req
      -- 
    req_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(370), ack => WPIPE_input_pipe4_506_inst_req_0); -- 
    access_T_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(100) & access_T_CP_0_elements(197) & access_T_CP_0_elements(235) & access_T_CP_0_elements(372);
      gj_access_T_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	96 
    -- CP-element group 371: 	193 
    -- CP-element group 371: 	231 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_update_start_
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Sample/ack
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Update/req
      -- 
    ack_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_506_inst_ack_0, ack => access_T_CP_0_elements(371)); -- 
    req_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(371), ack => WPIPE_input_pipe4_506_inst_req_1); -- 
    -- CP-element group 372:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: marked-successors 
    -- CP-element group 372: 	370 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/WPIPE_input_pipe4_506_Update/ack
      -- 
    ack_1590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_506_inst_ack_1, ack => access_T_CP_0_elements(372)); -- 
    -- CP-element group 373:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	30 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	31 
    -- CP-element group 373:  members (1) 
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(373) is a control-delay.
    cp_element_373_delay: control_delay_element  generic map(name => " 373_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(30), ack => access_T_CP_0_elements(373), clk => clk, reset =>reset);
    -- CP-element group 374:  join  transition  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	33 
    -- CP-element group 374: 	257 
    -- CP-element group 374: 	268 
    -- CP-element group 374: 	272 
    -- CP-element group 374: 	276 
    -- CP-element group 374: 	285 
    -- CP-element group 374: 	296 
    -- CP-element group 374: 	300 
    -- CP-element group 374: 	304 
    -- CP-element group 374: 	313 
    -- CP-element group 374: 	324 
    -- CP-element group 374: 	328 
    -- CP-element group 374: 	332 
    -- CP-element group 374: 	341 
    -- CP-element group 374: 	352 
    -- CP-element group 374: 	356 
    -- CP-element group 374: 	360 
    -- CP-element group 374: 	363 
    -- CP-element group 374: 	366 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	27 
    -- CP-element group 374:  members (1) 
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_100/do_while_stmt_100_loop_body/$exit
      -- 
    access_T_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15,20 => 15);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= access_T_CP_0_elements(33) & access_T_CP_0_elements(257) & access_T_CP_0_elements(268) & access_T_CP_0_elements(272) & access_T_CP_0_elements(276) & access_T_CP_0_elements(285) & access_T_CP_0_elements(296) & access_T_CP_0_elements(300) & access_T_CP_0_elements(304) & access_T_CP_0_elements(313) & access_T_CP_0_elements(324) & access_T_CP_0_elements(328) & access_T_CP_0_elements(332) & access_T_CP_0_elements(341) & access_T_CP_0_elements(352) & access_T_CP_0_elements(356) & access_T_CP_0_elements(360) & access_T_CP_0_elements(363) & access_T_CP_0_elements(366) & access_T_CP_0_elements(369) & access_T_CP_0_elements(372);
      gj_access_T_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	26 
    -- CP-element group 375: successors 
    -- CP-element group 375:  members (2) 
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_100/loop_exit/$exit
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_100/loop_exit/ack
      -- 
    ack_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_100_branch_ack_0, ack => access_T_CP_0_elements(375)); -- 
    -- CP-element group 376:  transition  input  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	26 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (2) 
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_100/loop_taken/$exit
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_100/loop_taken/ack
      -- 
    ack_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_100_branch_ack_1, ack => access_T_CP_0_elements(376)); -- 
    -- CP-element group 377:  transition  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	24 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	1 
    -- CP-element group 377:  members (1) 
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_100/$exit
      -- 
    access_T_CP_0_elements(377) <= access_T_CP_0_elements(24);
    access_T_do_while_stmt_100_terminator_1600: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_100_terminator_1600", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(27),loop_continue => access_T_CP_0_elements(376),loop_terminate => access_T_CP_0_elements(375),loop_back => access_T_CP_0_elements(25),loop_exit => access_T_CP_0_elements(24),clk => clk, reset => reset); -- 
    phi_stmt_102_phi_seq_416_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(44);
      access_T_CP_0_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(49);
      access_T_CP_0_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(53);
      access_T_CP_0_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(54);
      access_T_CP_0_elements(43) <= phi_mux_reqs(1);
      phi_stmt_102_phi_seq_416 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_102_phi_seq_416") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(38), 
          phi_sample_ack => access_T_CP_0_elements(39), 
          phi_update_req => access_T_CP_0_elements(40), 
          phi_update_ack => access_T_CP_0_elements(41), 
          phi_mux_ack => access_T_CP_0_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_107_phi_seq_470_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(63);
      access_T_CP_0_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(70);
      access_T_CP_0_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(71);
      access_T_CP_0_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(61);
      access_T_CP_0_elements(72)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(74);
      access_T_CP_0_elements(73)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(75);
      access_T_CP_0_elements(62) <= phi_mux_reqs(1);
      phi_stmt_107_phi_seq_470 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_107_phi_seq_470") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(57), 
          phi_sample_ack => access_T_CP_0_elements(58), 
          phi_update_req => access_T_CP_0_elements(59), 
          phi_update_ack => access_T_CP_0_elements(60), 
          phi_mux_ack => access_T_CP_0_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_112_phi_seq_524_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(82);
      access_T_CP_0_elements(85)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(89);
      access_T_CP_0_elements(86)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(90);
      access_T_CP_0_elements(83) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(80);
      access_T_CP_0_elements(91)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(93);
      access_T_CP_0_elements(92)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(94);
      access_T_CP_0_elements(81) <= phi_mux_reqs(1);
      phi_stmt_112_phi_seq_524 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_112_phi_seq_524") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(32), 
          phi_sample_ack => access_T_CP_0_elements(78), 
          phi_update_req => access_T_CP_0_elements(34), 
          phi_update_ack => access_T_CP_0_elements(79), 
          phi_mux_ack => access_T_CP_0_elements(84), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_117_phi_seq_578_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(103);
      access_T_CP_0_elements(106)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(110);
      access_T_CP_0_elements(107)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(111);
      access_T_CP_0_elements(104) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(101);
      access_T_CP_0_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(114);
      access_T_CP_0_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(115);
      access_T_CP_0_elements(102) <= phi_mux_reqs(1);
      phi_stmt_117_phi_seq_578 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_117_phi_seq_578") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(97), 
          phi_sample_ack => access_T_CP_0_elements(98), 
          phi_update_req => access_T_CP_0_elements(99), 
          phi_update_ack => access_T_CP_0_elements(100), 
          phi_mux_ack => access_T_CP_0_elements(105), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_124_phi_seq_622_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(124);
      access_T_CP_0_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(129);
      access_T_CP_0_elements(125) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(122);
      access_T_CP_0_elements(131)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(133);
      access_T_CP_0_elements(132)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(134);
      access_T_CP_0_elements(123) <= phi_mux_reqs(1);
      phi_stmt_124_phi_seq_622 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_124_phi_seq_622") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(118), 
          phi_sample_ack => access_T_CP_0_elements(119), 
          phi_update_req => access_T_CP_0_elements(120), 
          phi_update_ack => access_T_CP_0_elements(121), 
          phi_mux_ack => access_T_CP_0_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_129_phi_seq_676_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(143);
      access_T_CP_0_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(148);
      access_T_CP_0_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(149);
      access_T_CP_0_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(141);
      access_T_CP_0_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(152);
      access_T_CP_0_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(153);
      access_T_CP_0_elements(142) <= phi_mux_reqs(1);
      phi_stmt_129_phi_seq_676 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_129_phi_seq_676") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(137), 
          phi_sample_ack => access_T_CP_0_elements(138), 
          phi_update_req => access_T_CP_0_elements(139), 
          phi_update_ack => access_T_CP_0_elements(140), 
          phi_mux_ack => access_T_CP_0_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_133_phi_seq_730_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(162);
      access_T_CP_0_elements(165)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(167);
      access_T_CP_0_elements(166)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(168);
      access_T_CP_0_elements(163) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(160);
      access_T_CP_0_elements(169)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(171);
      access_T_CP_0_elements(170)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(172);
      access_T_CP_0_elements(161) <= phi_mux_reqs(1);
      phi_stmt_133_phi_seq_730 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_133_phi_seq_730") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(156), 
          phi_sample_ack => access_T_CP_0_elements(157), 
          phi_update_req => access_T_CP_0_elements(158), 
          phi_update_ack => access_T_CP_0_elements(159), 
          phi_mux_ack => access_T_CP_0_elements(164), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_137_phi_seq_784_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(181);
      access_T_CP_0_elements(184)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(186);
      access_T_CP_0_elements(185)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(187);
      access_T_CP_0_elements(182) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(179);
      access_T_CP_0_elements(188)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(190);
      access_T_CP_0_elements(189)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(191);
      access_T_CP_0_elements(180) <= phi_mux_reqs(1);
      phi_stmt_137_phi_seq_784 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_137_phi_seq_784") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(175), 
          phi_sample_ack => access_T_CP_0_elements(176), 
          phi_update_req => access_T_CP_0_elements(177), 
          phi_update_ack => access_T_CP_0_elements(178), 
          phi_mux_ack => access_T_CP_0_elements(183), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_141_phi_seq_838_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(200);
      access_T_CP_0_elements(203)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(205);
      access_T_CP_0_elements(204)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(206);
      access_T_CP_0_elements(201) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(198);
      access_T_CP_0_elements(207)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(209);
      access_T_CP_0_elements(208)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(210);
      access_T_CP_0_elements(199) <= phi_mux_reqs(1);
      phi_stmt_141_phi_seq_838 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_141_phi_seq_838") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(194), 
          phi_sample_ack => access_T_CP_0_elements(195), 
          phi_update_req => access_T_CP_0_elements(196), 
          phi_update_ack => access_T_CP_0_elements(197), 
          phi_mux_ack => access_T_CP_0_elements(202), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_145_phi_seq_882_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(219);
      access_T_CP_0_elements(222)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(222);
      access_T_CP_0_elements(223)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(224);
      access_T_CP_0_elements(220) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(217);
      access_T_CP_0_elements(226)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(228);
      access_T_CP_0_elements(227)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(229);
      access_T_CP_0_elements(218) <= phi_mux_reqs(1);
      phi_stmt_145_phi_seq_882 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_145_phi_seq_882") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(213), 
          phi_sample_ack => access_T_CP_0_elements(214), 
          phi_update_req => access_T_CP_0_elements(215), 
          phi_update_ack => access_T_CP_0_elements(216), 
          phi_mux_ack => access_T_CP_0_elements(221), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_150_phi_seq_926_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(238);
      access_T_CP_0_elements(241)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(241);
      access_T_CP_0_elements(242)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(243);
      access_T_CP_0_elements(239) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(236);
      access_T_CP_0_elements(245)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(247);
      access_T_CP_0_elements(246)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(248);
      access_T_CP_0_elements(237) <= phi_mux_reqs(1);
      phi_stmt_150_phi_seq_926 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_150_phi_seq_926") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(232), 
          phi_sample_ack => access_T_CP_0_elements(233), 
          phi_update_req => access_T_CP_0_elements(234), 
          phi_update_ack => access_T_CP_0_elements(235), 
          phi_mux_ack => access_T_CP_0_elements(240), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_368_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(28);
        preds(1)  <= access_T_CP_0_elements(29);
        entry_tmerge_368 : transition_merge -- 
          generic map(name => " entry_tmerge_368")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(30));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_183_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_191_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_121_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_166_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_91_wire : std_logic_vector(31 downto 0);
    signal ADD_u64_u64_233_wire : std_logic_vector(63 downto 0);
    signal ADD_u64_u64_305_wire : std_logic_vector(63 downto 0);
    signal ADD_u64_u64_377_wire : std_logic_vector(63 downto 0);
    signal ADD_u64_u64_449_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_209_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_281_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_353_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_425_wire : std_logic_vector(63 downto 0);
    signal LSHR_u32_u32_59_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_73_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_87_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_90_wire : std_logic_vector(31 downto 0);
    signal LSHR_u64_u64_217_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_240_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_243_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_253_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_253_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_253_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_289_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_312_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_315_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_325_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_325_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_325_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_361_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_384_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_387_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_397_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_397_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_397_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_433_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_456_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_459_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_469_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_469_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_469_wire : std_logic_vector(63 downto 0);
    signal MUL_u16_u16_34_wire : std_logic_vector(15 downto 0);
    signal NEQ_u64_u1_244_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_316_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_388_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_460_wire : std_logic_vector(0 downto 0);
    signal SUB_u64_u64_210_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_282_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_354_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_426_wire : std_logic_vector(63 downto 0);
    signal address1_102 : std_logic_vector(63 downto 0);
    signal address2_107 : std_logic_vector(63 downto 0);
    signal address3_112 : std_logic_vector(63 downto 0);
    signal address4_117 : std_logic_vector(63 downto 0);
    signal array_obj_ref_254_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_254_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_326_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_398_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_470_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_61_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_75_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_93_root_address : std_logic_vector(13 downto 0);
    signal continue1_199 : std_logic_vector(0 downto 0);
    signal continue2_204 : std_logic_vector(0 downto 0);
    signal fetch_add1_49 : std_logic_vector(31 downto 0);
    signal fetch_add2_63 : std_logic_vector(31 downto 0);
    signal fetch_add3_77 : std_logic_vector(31 downto 0);
    signal fetch_add4_95 : std_logic_vector(31 downto 0);
    signal fetch_addr1_256 : std_logic_vector(31 downto 0);
    signal fetch_addr2_328 : std_logic_vector(31 downto 0);
    signal fetch_addr3_400 : std_logic_vector(31 downto 0);
    signal fetch_addr4_472 : std_logic_vector(31 downto 0);
    signal fetch_val1_129 : std_logic_vector(63 downto 0);
    signal fetch_val1_262_delayed_13_0_270 : std_logic_vector(63 downto 0);
    signal fetch_val2_133 : std_logic_vector(63 downto 0);
    signal fetch_val2_322_delayed_13_0_342 : std_logic_vector(63 downto 0);
    signal fetch_val3_137 : std_logic_vector(63 downto 0);
    signal fetch_val3_382_delayed_13_0_414 : std_logic_vector(63 downto 0);
    signal fetch_val4_141 : std_logic_vector(63 downto 0);
    signal fetch_val4_442_delayed_13_0_486 : std_logic_vector(63 downto 0);
    signal fn1_247 : std_logic_vector(0 downto 0);
    signal fn1_254_delayed_7_0_259 : std_logic_vector(0 downto 0);
    signal fn1_260_delayed_13_0_267 : std_logic_vector(0 downto 0);
    signal fn2_314_delayed_7_0_331 : std_logic_vector(0 downto 0);
    signal fn2_319 : std_logic_vector(0 downto 0);
    signal fn2_320_delayed_13_0_339 : std_logic_vector(0 downto 0);
    signal fn3_374_delayed_7_0_403 : std_logic_vector(0 downto 0);
    signal fn3_380_delayed_13_0_411 : std_logic_vector(0 downto 0);
    signal fn3_391 : std_logic_vector(0 downto 0);
    signal fn4_434_delayed_7_0_475 : std_logic_vector(0 downto 0);
    signal fn4_440_delayed_13_0_483 : std_logic_vector(0 downto 0);
    signal fn4_463 : std_logic_vector(0 downto 0);
    signal fv1_264 : std_logic_vector(63 downto 0);
    signal fv2_336 : std_logic_vector(63 downto 0);
    signal fv3_408 : std_logic_vector(63 downto 0);
    signal fv4_480 : std_logic_vector(63 downto 0);
    signal konst_163_wire_constant : std_logic_vector(31 downto 0);
    signal konst_165_wire_constant : std_logic_vector(31 downto 0);
    signal konst_182_wire_constant : std_logic_vector(15 downto 0);
    signal konst_190_wire_constant : std_logic_vector(15 downto 0);
    signal konst_206_wire_constant : std_logic_vector(63 downto 0);
    signal konst_208_wire_constant : std_logic_vector(63 downto 0);
    signal konst_211_wire_constant : std_logic_vector(63 downto 0);
    signal konst_222_wire_constant : std_logic_vector(63 downto 0);
    signal konst_239_wire_constant : std_logic_vector(63 downto 0);
    signal konst_242_wire_constant : std_logic_vector(63 downto 0);
    signal konst_252_wire_constant : std_logic_vector(63 downto 0);
    signal konst_278_wire_constant : std_logic_vector(63 downto 0);
    signal konst_280_wire_constant : std_logic_vector(63 downto 0);
    signal konst_283_wire_constant : std_logic_vector(63 downto 0);
    signal konst_294_wire_constant : std_logic_vector(63 downto 0);
    signal konst_311_wire_constant : std_logic_vector(63 downto 0);
    signal konst_314_wire_constant : std_logic_vector(63 downto 0);
    signal konst_324_wire_constant : std_logic_vector(63 downto 0);
    signal konst_350_wire_constant : std_logic_vector(63 downto 0);
    signal konst_352_wire_constant : std_logic_vector(63 downto 0);
    signal konst_355_wire_constant : std_logic_vector(63 downto 0);
    signal konst_366_wire_constant : std_logic_vector(63 downto 0);
    signal konst_383_wire_constant : std_logic_vector(63 downto 0);
    signal konst_386_wire_constant : std_logic_vector(63 downto 0);
    signal konst_396_wire_constant : std_logic_vector(63 downto 0);
    signal konst_39_wire_constant : std_logic_vector(31 downto 0);
    signal konst_422_wire_constant : std_logic_vector(63 downto 0);
    signal konst_424_wire_constant : std_logic_vector(63 downto 0);
    signal konst_427_wire_constant : std_logic_vector(63 downto 0);
    signal konst_438_wire_constant : std_logic_vector(63 downto 0);
    signal konst_455_wire_constant : std_logic_vector(63 downto 0);
    signal konst_458_wire_constant : std_logic_vector(63 downto 0);
    signal konst_468_wire_constant : std_logic_vector(63 downto 0);
    signal konst_58_wire_constant : std_logic_vector(31 downto 0);
    signal konst_72_wire_constant : std_logic_vector(31 downto 0);
    signal konst_86_wire_constant : std_logic_vector(31 downto 0);
    signal konst_89_wire_constant : std_logic_vector(31 downto 0);
    signal m2_factor_41 : std_logic_vector(31 downto 0);
    signal m_factor_36 : std_logic_vector(31 downto 0);
    signal my_fetch1_53 : std_logic_vector(63 downto 0);
    signal my_fetch1_53_131_buffered : std_logic_vector(63 downto 0);
    signal my_fetch2_67 : std_logic_vector(63 downto 0);
    signal my_fetch2_67_135_buffered : std_logic_vector(63 downto 0);
    signal my_fetch3_81 : std_logic_vector(63 downto 0);
    signal my_fetch3_81_139_buffered : std_logic_vector(63 downto 0);
    signal my_fetch4_99 : std_logic_vector(63 downto 0);
    signal my_fetch4_99_143_buffered : std_logic_vector(63 downto 0);
    signal my_num1_213 : std_logic_vector(63 downto 0);
    signal my_num2_285 : std_logic_vector(63 downto 0);
    signal my_num3_357 : std_logic_vector(63 downto 0);
    signal my_num4_429 : std_logic_vector(63 downto 0);
    signal mycounter_124 : std_logic_vector(31 downto 0);
    signal n_address1_236 : std_logic_vector(63 downto 0);
    signal n_address1_236_106_buffered : std_logic_vector(63 downto 0);
    signal n_address2_308 : std_logic_vector(63 downto 0);
    signal n_address2_308_111_buffered : std_logic_vector(63 downto 0);
    signal n_address3_380 : std_logic_vector(63 downto 0);
    signal n_address3_380_116_buffered : std_logic_vector(63 downto 0);
    signal n_address4_452 : std_logic_vector(63 downto 0);
    signal n_address4_452_123_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val1_276 : std_logic_vector(63 downto 0);
    signal n_fetch_val1_276_132_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val2_348 : std_logic_vector(63 downto 0);
    signal n_fetch_val2_348_136_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val3_420 : std_logic_vector(63 downto 0);
    signal n_fetch_val3_420_140_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val4_492 : std_logic_vector(63 downto 0);
    signal n_fetch_val4_492_144_buffered : std_logic_vector(63 downto 0);
    signal n_mycounter_168 : std_logic_vector(31 downto 0);
    signal n_mycounter_168_128_buffered : std_logic_vector(31 downto 0);
    signal n_row1_186 : std_logic_vector(15 downto 0);
    signal n_row1_186_149_buffered : std_logic_vector(15 downto 0);
    signal n_row2_194 : std_logic_vector(15 downto 0);
    signal n_row2_194_154_buffered : std_logic_vector(15 downto 0);
    signal next_row_160 : std_logic_vector(0 downto 0);
    signal ptr_deref_263_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_263_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_263_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_263_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_263_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_335_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_335_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_335_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_335_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_335_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_407_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_407_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_407_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_407_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_407_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_479_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_479_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_479_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_479_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_479_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_52_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_52_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_52_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_52_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_52_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_66_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_66_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_66_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_66_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_66_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_80_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_80_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_80_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_80_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_80_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_98_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_98_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_98_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_98_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_98_word_offset_0 : std_logic_vector(13 downto 0);
    signal row1_145 : std_logic_vector(15 downto 0);
    signal row2_150 : std_logic_vector(15 downto 0);
    signal send_now1_173 : std_logic_vector(0 downto 0);
    signal send_now2_178 : std_logic_vector(0 downto 0);
    signal temp_address1_224 : std_logic_vector(63 downto 0);
    signal temp_address2_296 : std_logic_vector(63 downto 0);
    signal temp_address3_368 : std_logic_vector(63 downto 0);
    signal temp_address4_440 : std_logic_vector(63 downto 0);
    signal type_cast_105_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_110_wire : std_logic_vector(63 downto 0);
    signal type_cast_115_wire : std_logic_vector(63 downto 0);
    signal type_cast_122_wire : std_logic_vector(63 downto 0);
    signal type_cast_127_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_148_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_153_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_229_229_delayed_1_0_228 : std_logic_vector(63 downto 0);
    signal type_cast_289_289_delayed_1_0_300 : std_logic_vector(63 downto 0);
    signal type_cast_349_349_delayed_1_0_372 : std_logic_vector(63 downto 0);
    signal type_cast_409_409_delayed_1_0_444 : std_logic_vector(63 downto 0);
    signal type_cast_60_resized : std_logic_vector(13 downto 0);
    signal type_cast_60_scaled : std_logic_vector(13 downto 0);
    signal type_cast_60_wire : std_logic_vector(63 downto 0);
    signal type_cast_74_resized : std_logic_vector(13 downto 0);
    signal type_cast_74_scaled : std_logic_vector(13 downto 0);
    signal type_cast_74_wire : std_logic_vector(63 downto 0);
    signal type_cast_92_resized : std_logic_vector(13 downto 0);
    signal type_cast_92_scaled : std_logic_vector(13 downto 0);
    signal type_cast_92_wire : std_logic_vector(63 downto 0);
    signal var_val1_219 : std_logic_vector(15 downto 0);
    signal var_val2_291 : std_logic_vector(15 downto 0);
    signal var_val3_363 : std_logic_vector(15 downto 0);
    signal var_val4_435 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_254_constant_part_of_offset <= "00000000000000";
    array_obj_ref_254_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_254_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_254_resized_base_address <= "00000000000000";
    array_obj_ref_326_constant_part_of_offset <= "00000000000000";
    array_obj_ref_326_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_326_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_326_resized_base_address <= "00000000000000";
    array_obj_ref_398_constant_part_of_offset <= "00000000000000";
    array_obj_ref_398_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_398_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_398_resized_base_address <= "00000000000000";
    array_obj_ref_470_constant_part_of_offset <= "00000000000000";
    array_obj_ref_470_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_470_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_470_resized_base_address <= "00000000000000";
    array_obj_ref_61_constant_part_of_offset <= "00000000000000";
    array_obj_ref_61_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_61_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_61_resized_base_address <= "00000000000000";
    array_obj_ref_75_constant_part_of_offset <= "00000000000000";
    array_obj_ref_75_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_75_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_75_resized_base_address <= "00000000000000";
    array_obj_ref_93_constant_part_of_offset <= "00000000000000";
    array_obj_ref_93_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_93_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_93_resized_base_address <= "00000000000000";
    fetch_add1_49 <= "00000000000000000000000000000000";
    konst_163_wire_constant <= "00000000000000000000000000000001";
    konst_165_wire_constant <= "00000000000000000000000000000001";
    konst_182_wire_constant <= "0000000000000010";
    konst_190_wire_constant <= "0000000000000010";
    konst_206_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_208_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_211_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_222_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_239_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_242_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_252_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_278_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_280_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_283_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_294_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_311_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_314_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_324_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_350_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_352_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_355_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_366_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_383_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_396_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_39_wire_constant <= "00000000000000000000000000000001";
    konst_422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_424_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_427_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_455_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_458_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_468_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_58_wire_constant <= "00000000000000000000000000000010";
    konst_72_wire_constant <= "00000000000000000000000000000001";
    konst_86_wire_constant <= "00000000000000000000000000000001";
    konst_89_wire_constant <= "00000000000000000000000000000010";
    ptr_deref_263_word_offset_0 <= "00000000000000";
    ptr_deref_335_word_offset_0 <= "00000000000000";
    ptr_deref_407_word_offset_0 <= "00000000000000";
    ptr_deref_479_word_offset_0 <= "00000000000000";
    ptr_deref_52_word_offset_0 <= "00000000000000";
    ptr_deref_66_word_offset_0 <= "00000000000000";
    ptr_deref_80_word_offset_0 <= "00000000000000";
    ptr_deref_98_word_offset_0 <= "00000000000000";
    type_cast_105_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_127_wire_constant <= "00000000000000000000000000000001";
    type_cast_148_wire_constant <= "0000000000000000";
    type_cast_153_wire_constant <= "0000000000000001";
    phi_stmt_102: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_105_wire_constant & n_address1_236_106_buffered;
      req <= phi_stmt_102_req_0 & phi_stmt_102_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_102",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_102_ack_0,
          idata => idata,
          odata => address1_102,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_102
    phi_stmt_107: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_110_wire & n_address2_308_111_buffered;
      req <= phi_stmt_107_req_0 & phi_stmt_107_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_107",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_107_ack_0,
          idata => idata,
          odata => address2_107,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_107
    phi_stmt_112: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_115_wire & n_address3_380_116_buffered;
      req <= phi_stmt_112_req_0 & phi_stmt_112_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_112",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_112_ack_0,
          idata => idata,
          odata => address3_112,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_112
    phi_stmt_117: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_122_wire & n_address4_452_123_buffered;
      req <= phi_stmt_117_req_0 & phi_stmt_117_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_117",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_117_ack_0,
          idata => idata,
          odata => address4_117,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_117
    phi_stmt_124: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_127_wire_constant & n_mycounter_168_128_buffered;
      req <= phi_stmt_124_req_0 & phi_stmt_124_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_124",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_124_ack_0,
          idata => idata,
          odata => mycounter_124,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_124
    phi_stmt_129: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch1_53_131_buffered & n_fetch_val1_276_132_buffered;
      req <= phi_stmt_129_req_0 & phi_stmt_129_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_129",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_129_ack_0,
          idata => idata,
          odata => fetch_val1_129,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_129
    phi_stmt_133: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch2_67_135_buffered & n_fetch_val2_348_136_buffered;
      req <= phi_stmt_133_req_0 & phi_stmt_133_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_133",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_133_ack_0,
          idata => idata,
          odata => fetch_val2_133,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_133
    phi_stmt_137: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch3_81_139_buffered & n_fetch_val3_420_140_buffered;
      req <= phi_stmt_137_req_0 & phi_stmt_137_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_137",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_137_ack_0,
          idata => idata,
          odata => fetch_val3_137,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_137
    phi_stmt_141: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch4_99_143_buffered & n_fetch_val4_492_144_buffered;
      req <= phi_stmt_141_req_0 & phi_stmt_141_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_141",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_141_ack_0,
          idata => idata,
          odata => fetch_val4_141,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_141
    phi_stmt_145: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_148_wire_constant & n_row1_186_149_buffered;
      req <= phi_stmt_145_req_0 & phi_stmt_145_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_145",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_145_ack_0,
          idata => idata,
          odata => row1_145,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_145
    phi_stmt_150: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_153_wire_constant & n_row2_194_154_buffered;
      req <= phi_stmt_150_req_0 & phi_stmt_150_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_150",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_150_ack_0,
          idata => idata,
          odata => row2_150,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_150
    -- flow-through select operator MUX_167_inst
    n_mycounter_168 <= konst_163_wire_constant when (next_row_160(0) /=  '0') else ADD_u32_u32_166_wire;
    -- flow-through select operator MUX_185_inst
    n_row1_186 <= ADD_u16_u16_183_wire when (next_row_160(0) /=  '0') else row1_145;
    -- flow-through select operator MUX_193_inst
    n_row2_194 <= ADD_u16_u16_191_wire when (next_row_160(0) /=  '0') else row2_150;
    -- flow-through select operator MUX_235_inst
    n_address1_236 <= ADD_u64_u64_233_wire when (next_row_160(0) /=  '0') else temp_address1_224;
    -- flow-through select operator MUX_275_inst
    n_fetch_val1_276 <= fv1_264 when (fn1_260_delayed_13_0_267(0) /=  '0') else fetch_val1_262_delayed_13_0_270;
    -- flow-through select operator MUX_307_inst
    n_address2_308 <= ADD_u64_u64_305_wire when (next_row_160(0) /=  '0') else temp_address2_296;
    -- flow-through select operator MUX_347_inst
    n_fetch_val2_348 <= fv2_336 when (fn2_320_delayed_13_0_339(0) /=  '0') else fetch_val2_322_delayed_13_0_342;
    -- flow-through select operator MUX_379_inst
    n_address3_380 <= ADD_u64_u64_377_wire when (next_row_160(0) /=  '0') else temp_address3_368;
    -- flow-through select operator MUX_419_inst
    n_fetch_val3_420 <= fv3_408 when (fn3_380_delayed_13_0_411(0) /=  '0') else fetch_val3_382_delayed_13_0_414;
    -- flow-through select operator MUX_451_inst
    n_address4_452 <= ADD_u64_u64_449_wire when (next_row_160(0) /=  '0') else temp_address4_440;
    -- flow-through select operator MUX_491_inst
    n_fetch_val4_492 <= fv4_480 when (fn4_440_delayed_13_0_483(0) /=  '0') else fetch_val4_442_delayed_13_0_486;
    W_fetch_val1_262_delayed_13_0_268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val1_262_delayed_13_0_268_inst_req_0;
      W_fetch_val1_262_delayed_13_0_268_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val1_262_delayed_13_0_268_inst_req_1;
      W_fetch_val1_262_delayed_13_0_268_inst_ack_1<= rack(0);
      W_fetch_val1_262_delayed_13_0_268_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val1_262_delayed_13_0_268_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val1_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val1_262_delayed_13_0_270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val2_322_delayed_13_0_340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val2_322_delayed_13_0_340_inst_req_0;
      W_fetch_val2_322_delayed_13_0_340_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val2_322_delayed_13_0_340_inst_req_1;
      W_fetch_val2_322_delayed_13_0_340_inst_ack_1<= rack(0);
      W_fetch_val2_322_delayed_13_0_340_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val2_322_delayed_13_0_340_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val2_133,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val2_322_delayed_13_0_342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val3_382_delayed_13_0_412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val3_382_delayed_13_0_412_inst_req_0;
      W_fetch_val3_382_delayed_13_0_412_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val3_382_delayed_13_0_412_inst_req_1;
      W_fetch_val3_382_delayed_13_0_412_inst_ack_1<= rack(0);
      W_fetch_val3_382_delayed_13_0_412_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val3_382_delayed_13_0_412_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val3_137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val3_382_delayed_13_0_414,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val4_442_delayed_13_0_484_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val4_442_delayed_13_0_484_inst_req_0;
      W_fetch_val4_442_delayed_13_0_484_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val4_442_delayed_13_0_484_inst_req_1;
      W_fetch_val4_442_delayed_13_0_484_inst_ack_1<= rack(0);
      W_fetch_val4_442_delayed_13_0_484_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val4_442_delayed_13_0_484_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val4_141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val4_442_delayed_13_0_486,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn1_254_delayed_7_0_257_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn1_254_delayed_7_0_257_inst_req_0;
      W_fn1_254_delayed_7_0_257_inst_ack_0<= wack(0);
      rreq(0) <= W_fn1_254_delayed_7_0_257_inst_req_1;
      W_fn1_254_delayed_7_0_257_inst_ack_1<= rack(0);
      W_fn1_254_delayed_7_0_257_inst : InterlockBuffer generic map ( -- 
        name => "W_fn1_254_delayed_7_0_257_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn1_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn1_254_delayed_7_0_259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn1_260_delayed_13_0_265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn1_260_delayed_13_0_265_inst_req_0;
      W_fn1_260_delayed_13_0_265_inst_ack_0<= wack(0);
      rreq(0) <= W_fn1_260_delayed_13_0_265_inst_req_1;
      W_fn1_260_delayed_13_0_265_inst_ack_1<= rack(0);
      W_fn1_260_delayed_13_0_265_inst : InterlockBuffer generic map ( -- 
        name => "W_fn1_260_delayed_13_0_265_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn1_247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn1_260_delayed_13_0_267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn2_314_delayed_7_0_329_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn2_314_delayed_7_0_329_inst_req_0;
      W_fn2_314_delayed_7_0_329_inst_ack_0<= wack(0);
      rreq(0) <= W_fn2_314_delayed_7_0_329_inst_req_1;
      W_fn2_314_delayed_7_0_329_inst_ack_1<= rack(0);
      W_fn2_314_delayed_7_0_329_inst : InterlockBuffer generic map ( -- 
        name => "W_fn2_314_delayed_7_0_329_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn2_319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn2_314_delayed_7_0_331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn2_320_delayed_13_0_337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn2_320_delayed_13_0_337_inst_req_0;
      W_fn2_320_delayed_13_0_337_inst_ack_0<= wack(0);
      rreq(0) <= W_fn2_320_delayed_13_0_337_inst_req_1;
      W_fn2_320_delayed_13_0_337_inst_ack_1<= rack(0);
      W_fn2_320_delayed_13_0_337_inst : InterlockBuffer generic map ( -- 
        name => "W_fn2_320_delayed_13_0_337_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn2_319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn2_320_delayed_13_0_339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn3_374_delayed_7_0_401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn3_374_delayed_7_0_401_inst_req_0;
      W_fn3_374_delayed_7_0_401_inst_ack_0<= wack(0);
      rreq(0) <= W_fn3_374_delayed_7_0_401_inst_req_1;
      W_fn3_374_delayed_7_0_401_inst_ack_1<= rack(0);
      W_fn3_374_delayed_7_0_401_inst : InterlockBuffer generic map ( -- 
        name => "W_fn3_374_delayed_7_0_401_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn3_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn3_374_delayed_7_0_403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn3_380_delayed_13_0_409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn3_380_delayed_13_0_409_inst_req_0;
      W_fn3_380_delayed_13_0_409_inst_ack_0<= wack(0);
      rreq(0) <= W_fn3_380_delayed_13_0_409_inst_req_1;
      W_fn3_380_delayed_13_0_409_inst_ack_1<= rack(0);
      W_fn3_380_delayed_13_0_409_inst : InterlockBuffer generic map ( -- 
        name => "W_fn3_380_delayed_13_0_409_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn3_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn3_380_delayed_13_0_411,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn4_434_delayed_7_0_473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn4_434_delayed_7_0_473_inst_req_0;
      W_fn4_434_delayed_7_0_473_inst_ack_0<= wack(0);
      rreq(0) <= W_fn4_434_delayed_7_0_473_inst_req_1;
      W_fn4_434_delayed_7_0_473_inst_ack_1<= rack(0);
      W_fn4_434_delayed_7_0_473_inst : InterlockBuffer generic map ( -- 
        name => "W_fn4_434_delayed_7_0_473_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn4_463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn4_434_delayed_7_0_475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn4_440_delayed_13_0_481_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn4_440_delayed_13_0_481_inst_req_0;
      W_fn4_440_delayed_13_0_481_inst_ack_0<= wack(0);
      rreq(0) <= W_fn4_440_delayed_13_0_481_inst_req_1;
      W_fn4_440_delayed_13_0_481_inst_ack_1<= rack(0);
      W_fn4_440_delayed_13_0_481_inst : InterlockBuffer generic map ( -- 
        name => "W_fn4_440_delayed_13_0_481_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn4_463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn4_440_delayed_13_0_483,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_255_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_255_final_reg_req_0;
      addr_of_255_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_255_final_reg_req_1;
      addr_of_255_final_reg_ack_1<= rack(0);
      addr_of_255_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_255_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_254_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_327_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_327_final_reg_req_0;
      addr_of_327_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_327_final_reg_req_1;
      addr_of_327_final_reg_ack_1<= rack(0);
      addr_of_327_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_327_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_326_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_328,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_399_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_399_final_reg_req_0;
      addr_of_399_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_399_final_reg_req_1;
      addr_of_399_final_reg_ack_1<= rack(0);
      addr_of_399_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_399_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_398_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr3_400,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_471_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_471_final_reg_req_0;
      addr_of_471_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_471_final_reg_req_1;
      addr_of_471_final_reg_ack_1<= rack(0);
      addr_of_471_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_471_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_470_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr4_472,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_62_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_62_final_reg_req_0;
      addr_of_62_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_62_final_reg_req_1;
      addr_of_62_final_reg_ack_1<= rack(0);
      addr_of_62_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_62_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_61_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add2_63,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_76_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_76_final_reg_req_0;
      addr_of_76_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_76_final_reg_req_1;
      addr_of_76_final_reg_ack_1<= rack(0);
      addr_of_76_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_76_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_75_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add3_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_94_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_94_final_reg_req_0;
      addr_of_94_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_94_final_reg_req_1;
      addr_of_94_final_reg_ack_1<= rack(0);
      addr_of_94_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_94_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_93_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add4_95,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch1_53_131_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch1_53_131_buf_req_0;
      my_fetch1_53_131_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch1_53_131_buf_req_1;
      my_fetch1_53_131_buf_ack_1<= rack(0);
      my_fetch1_53_131_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch1_53_131_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch1_53,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch1_53_131_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch2_67_135_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch2_67_135_buf_req_0;
      my_fetch2_67_135_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch2_67_135_buf_req_1;
      my_fetch2_67_135_buf_ack_1<= rack(0);
      my_fetch2_67_135_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch2_67_135_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch2_67,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch2_67_135_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch3_81_139_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch3_81_139_buf_req_0;
      my_fetch3_81_139_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch3_81_139_buf_req_1;
      my_fetch3_81_139_buf_ack_1<= rack(0);
      my_fetch3_81_139_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch3_81_139_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch3_81,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch3_81_139_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch4_99_143_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch4_99_143_buf_req_0;
      my_fetch4_99_143_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch4_99_143_buf_req_1;
      my_fetch4_99_143_buf_ack_1<= rack(0);
      my_fetch4_99_143_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch4_99_143_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch4_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch4_99_143_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_236_106_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_236_106_buf_req_0;
      n_address1_236_106_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_236_106_buf_req_1;
      n_address1_236_106_buf_ack_1<= rack(0);
      n_address1_236_106_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_236_106_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_236,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_236_106_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_308_111_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_308_111_buf_req_0;
      n_address2_308_111_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_308_111_buf_req_1;
      n_address2_308_111_buf_ack_1<= rack(0);
      n_address2_308_111_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_308_111_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_308_111_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address3_380_116_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address3_380_116_buf_req_0;
      n_address3_380_116_buf_ack_0<= wack(0);
      rreq(0) <= n_address3_380_116_buf_req_1;
      n_address3_380_116_buf_ack_1<= rack(0);
      n_address3_380_116_buf : InterlockBuffer generic map ( -- 
        name => "n_address3_380_116_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address3_380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address3_380_116_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address4_452_123_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address4_452_123_buf_req_0;
      n_address4_452_123_buf_ack_0<= wack(0);
      rreq(0) <= n_address4_452_123_buf_req_1;
      n_address4_452_123_buf_ack_1<= rack(0);
      n_address4_452_123_buf : InterlockBuffer generic map ( -- 
        name => "n_address4_452_123_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address4_452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address4_452_123_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val1_276_132_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val1_276_132_buf_req_0;
      n_fetch_val1_276_132_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val1_276_132_buf_req_1;
      n_fetch_val1_276_132_buf_ack_1<= rack(0);
      n_fetch_val1_276_132_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val1_276_132_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val1_276,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val1_276_132_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val2_348_136_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val2_348_136_buf_req_0;
      n_fetch_val2_348_136_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val2_348_136_buf_req_1;
      n_fetch_val2_348_136_buf_ack_1<= rack(0);
      n_fetch_val2_348_136_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val2_348_136_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val2_348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val2_348_136_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val3_420_140_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val3_420_140_buf_req_0;
      n_fetch_val3_420_140_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val3_420_140_buf_req_1;
      n_fetch_val3_420_140_buf_ack_1<= rack(0);
      n_fetch_val3_420_140_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val3_420_140_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val3_420,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val3_420_140_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val4_492_144_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val4_492_144_buf_req_0;
      n_fetch_val4_492_144_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val4_492_144_buf_req_1;
      n_fetch_val4_492_144_buf_ack_1<= rack(0);
      n_fetch_val4_492_144_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val4_492_144_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val4_492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val4_492_144_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter_168_128_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter_168_128_buf_req_0;
      n_mycounter_168_128_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter_168_128_buf_req_1;
      n_mycounter_168_128_buf_ack_1<= rack(0);
      n_mycounter_168_128_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter_168_128_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter_168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter_168_128_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row1_186_149_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row1_186_149_buf_req_0;
      n_row1_186_149_buf_ack_0<= wack(0);
      rreq(0) <= n_row1_186_149_buf_req_1;
      n_row1_186_149_buf_ack_1<= rack(0);
      n_row1_186_149_buf : InterlockBuffer generic map ( -- 
        name => "n_row1_186_149_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row1_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row1_186_149_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row2_194_154_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row2_194_154_buf_req_0;
      n_row2_194_154_buf_ack_0<= wack(0);
      rreq(0) <= n_row2_194_154_buf_req_1;
      n_row2_194_154_buf_ack_1<= rack(0);
      n_row2_194_154_buf : InterlockBuffer generic map ( -- 
        name => "n_row2_194_154_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row2_194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row2_194_154_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_110_inst_req_0;
      type_cast_110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_110_inst_req_1;
      type_cast_110_inst_ack_1<= rack(0);
      type_cast_110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_110_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_110_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_115_inst_req_0;
      type_cast_115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_115_inst_req_1;
      type_cast_115_inst_ack_1<= rack(0);
      type_cast_115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_115_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m2_factor_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_115_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_122_inst_req_0;
      type_cast_122_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_122_inst_req_1;
      type_cast_122_inst_ack_1<= rack(0);
      type_cast_122_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_122_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u32_u32_121_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_122_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_218_inst
    process(LSHR_u64_u64_217_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_217_wire(15 downto 0);
      var_val1_219 <= tmp_var; -- 
    end process;
    type_cast_227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_227_inst_req_0;
      type_cast_227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_227_inst_req_1;
      type_cast_227_inst_ack_1<= rack(0);
      type_cast_227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_227_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_229_229_delayed_1_0_228,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_290_inst
    process(LSHR_u64_u64_289_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_289_wire(15 downto 0);
      var_val2_291 <= tmp_var; -- 
    end process;
    type_cast_299_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_299_inst_req_0;
      type_cast_299_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_299_inst_req_1;
      type_cast_299_inst_ack_1<= rack(0);
      type_cast_299_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_299_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_289_289_delayed_1_0_300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_35_inst
    process(MUL_u16_u16_34_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_34_wire(15 downto 0);
      m_factor_36 <= tmp_var; -- 
    end process;
    -- interlock type_cast_362_inst
    process(LSHR_u64_u64_361_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_361_wire(15 downto 0);
      var_val3_363 <= tmp_var; -- 
    end process;
    type_cast_371_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_371_inst_req_0;
      type_cast_371_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_371_inst_req_1;
      type_cast_371_inst_ack_1<= rack(0);
      type_cast_371_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_371_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_349_349_delayed_1_0_372,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_434_inst
    process(LSHR_u64_u64_433_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_433_wire(15 downto 0);
      var_val4_435 <= tmp_var; -- 
    end process;
    type_cast_443_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_443_inst_req_0;
      type_cast_443_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_443_inst_req_1;
      type_cast_443_inst_ack_1<= rack(0);
      type_cast_443_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_443_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_409_409_delayed_1_0_444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_60_inst
    process(LSHR_u32_u32_59_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_59_wire(31 downto 0);
      type_cast_60_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_74_inst
    process(LSHR_u32_u32_73_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_73_wire(31 downto 0);
      type_cast_74_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_92_inst
    process(ADD_u32_u32_91_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ADD_u32_u32_91_wire(31 downto 0);
      type_cast_92_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_254_index_1_rename
    process(LSHR_u64_u64_253_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_253_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_253_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_254_index_1_resize
    process(LSHR_u64_u64_253_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_253_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_253_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_254_root_address_inst
    process(array_obj_ref_254_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_254_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_254_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_326_index_1_rename
    process(LSHR_u64_u64_325_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_325_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_325_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_326_index_1_resize
    process(LSHR_u64_u64_325_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_325_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_325_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_326_root_address_inst
    process(array_obj_ref_326_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_326_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_326_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_index_1_rename
    process(LSHR_u64_u64_397_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_397_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_397_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_index_1_resize
    process(LSHR_u64_u64_397_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_397_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_397_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_root_address_inst
    process(array_obj_ref_398_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_398_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_398_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_470_index_1_rename
    process(LSHR_u64_u64_469_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_469_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_469_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_470_index_1_resize
    process(LSHR_u64_u64_469_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_469_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_469_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_470_root_address_inst
    process(array_obj_ref_470_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_470_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_470_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_index_1_rename
    process(type_cast_60_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_60_resized;
      ov(13 downto 0) := iv;
      type_cast_60_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_index_1_resize
    process(type_cast_60_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_60_wire;
      ov := iv(13 downto 0);
      type_cast_60_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_61_root_address_inst
    process(array_obj_ref_61_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_61_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_61_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_index_1_rename
    process(type_cast_74_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_74_resized;
      ov(13 downto 0) := iv;
      type_cast_74_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_index_1_resize
    process(type_cast_74_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_74_wire;
      ov := iv(13 downto 0);
      type_cast_74_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_75_root_address_inst
    process(array_obj_ref_75_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_75_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_75_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_index_1_rename
    process(type_cast_92_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_92_resized;
      ov(13 downto 0) := iv;
      type_cast_92_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_index_1_resize
    process(type_cast_92_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_92_wire;
      ov := iv(13 downto 0);
      type_cast_92_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_93_root_address_inst
    process(array_obj_ref_93_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_93_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_93_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_addr_0
    process(ptr_deref_263_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_263_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_263_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_base_resize
    process(fetch_addr1_256) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_256;
      ov := iv(13 downto 0);
      ptr_deref_263_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_gather_scatter
    process(ptr_deref_263_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_263_data_0;
      ov(63 downto 0) := iv;
      fv1_264 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_263_root_address_inst
    process(ptr_deref_263_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_263_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_263_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_335_addr_0
    process(ptr_deref_335_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_335_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_335_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_335_base_resize
    process(fetch_addr2_328) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_328;
      ov := iv(13 downto 0);
      ptr_deref_335_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_335_gather_scatter
    process(ptr_deref_335_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_335_data_0;
      ov(63 downto 0) := iv;
      fv2_336 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_335_root_address_inst
    process(ptr_deref_335_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_335_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_335_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_addr_0
    process(ptr_deref_407_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_407_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_base_resize
    process(fetch_addr3_400) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr3_400;
      ov := iv(13 downto 0);
      ptr_deref_407_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_gather_scatter
    process(ptr_deref_407_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_data_0;
      ov(63 downto 0) := iv;
      fv3_408 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_407_root_address_inst
    process(ptr_deref_407_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_407_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_407_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_addr_0
    process(ptr_deref_479_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_479_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_479_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_base_resize
    process(fetch_addr4_472) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr4_472;
      ov := iv(13 downto 0);
      ptr_deref_479_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_gather_scatter
    process(ptr_deref_479_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_479_data_0;
      ov(63 downto 0) := iv;
      fv4_480 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_479_root_address_inst
    process(ptr_deref_479_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_479_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_479_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_52_addr_0
    process(ptr_deref_52_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_52_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_52_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_52_base_resize
    process(fetch_add1_49) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add1_49;
      ov := iv(13 downto 0);
      ptr_deref_52_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_52_gather_scatter
    process(ptr_deref_52_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_52_data_0;
      ov(63 downto 0) := iv;
      my_fetch1_53 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_52_root_address_inst
    process(ptr_deref_52_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_52_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_52_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_addr_0
    process(ptr_deref_66_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_66_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_base_resize
    process(fetch_add2_63) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add2_63;
      ov := iv(13 downto 0);
      ptr_deref_66_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_gather_scatter
    process(ptr_deref_66_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_data_0;
      ov(63 downto 0) := iv;
      my_fetch2_67 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_root_address_inst
    process(ptr_deref_66_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_66_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_80_addr_0
    process(ptr_deref_80_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_80_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_80_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_80_base_resize
    process(fetch_add3_77) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add3_77;
      ov := iv(13 downto 0);
      ptr_deref_80_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_80_gather_scatter
    process(ptr_deref_80_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_80_data_0;
      ov(63 downto 0) := iv;
      my_fetch3_81 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_80_root_address_inst
    process(ptr_deref_80_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_80_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_80_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_98_addr_0
    process(ptr_deref_98_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_98_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_98_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_98_base_resize
    process(fetch_add4_95) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add4_95;
      ov := iv(13 downto 0);
      ptr_deref_98_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_98_gather_scatter
    process(ptr_deref_98_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_98_data_0;
      ov(63 downto 0) := iv;
      my_fetch4_99 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_98_root_address_inst
    process(ptr_deref_98_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_98_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_98_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_100_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue1_199;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_100_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_100_branch_req_0,
          ack0 => do_while_stmt_100_branch_ack_0,
          ack1 => do_while_stmt_100_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_183_inst
    process(row1_145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row1_145, konst_182_wire_constant, tmp_var);
      ADD_u16_u16_183_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_191_inst
    process(row2_150) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row2_150, konst_190_wire_constant, tmp_var);
      ADD_u16_u16_191_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_121_inst
    process(m_factor_36, m2_factor_41) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, m2_factor_41, tmp_var);
      ADD_u32_u32_121_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_166_inst
    process(mycounter_124) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycounter_124, konst_165_wire_constant, tmp_var);
      ADD_u32_u32_166_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_91_inst
    process(LSHR_u32_u32_87_wire, LSHR_u32_u32_90_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(LSHR_u32_u32_87_wire, LSHR_u32_u32_90_wire, tmp_var);
      ADD_u32_u32_91_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_223_inst
    process(address1_102) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_102, konst_222_wire_constant, tmp_var);
      temp_address1_224 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_233_inst
    process(temp_address1_224, type_cast_229_229_delayed_1_0_228) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(temp_address1_224, type_cast_229_229_delayed_1_0_228, tmp_var);
      ADD_u64_u64_233_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_295_inst
    process(address2_107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_107, konst_294_wire_constant, tmp_var);
      temp_address2_296 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_305_inst
    process(temp_address2_296, type_cast_289_289_delayed_1_0_300) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(temp_address2_296, type_cast_289_289_delayed_1_0_300, tmp_var);
      ADD_u64_u64_305_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_367_inst
    process(address3_112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address3_112, konst_366_wire_constant, tmp_var);
      temp_address3_368 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_377_inst
    process(temp_address3_368, type_cast_349_349_delayed_1_0_372) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(temp_address3_368, type_cast_349_349_delayed_1_0_372, tmp_var);
      ADD_u64_u64_377_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_439_inst
    process(address4_117) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address4_117, konst_438_wire_constant, tmp_var);
      temp_address4_440 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_449_inst
    process(temp_address4_440, type_cast_409_409_delayed_1_0_444) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(temp_address4_440, type_cast_409_409_delayed_1_0_444, tmp_var);
      ADD_u64_u64_449_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_246_inst
    process(NEQ_u64_u1_244_wire, continue1_199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_244_wire, continue1_199, tmp_var);
      fn1_247 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_318_inst
    process(NEQ_u64_u1_316_wire, continue1_199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_316_wire, continue1_199, tmp_var);
      fn2_319 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_390_inst
    process(NEQ_u64_u1_388_wire, continue1_199) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_388_wire, continue1_199, tmp_var);
      fn3_391 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_462_inst
    process(NEQ_u64_u1_460_wire, continue2_204) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_460_wire, continue2_204, tmp_var);
      fn4_463 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_209_inst
    process(address1_102) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address1_102, konst_208_wire_constant, tmp_var);
      AND_u64_u64_209_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_281_inst
    process(address2_107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address2_107, konst_280_wire_constant, tmp_var);
      AND_u64_u64_281_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_353_inst
    process(address3_112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address3_112, konst_352_wire_constant, tmp_var);
      AND_u64_u64_353_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_425_inst
    process(address4_117) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address4_117, konst_424_wire_constant, tmp_var);
      AND_u64_u64_425_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_159_inst
    process(mycounter_124, m_factor_36) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycounter_124, m_factor_36, tmp_var);
      next_row_160 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_59_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_36, konst_58_wire_constant, tmp_var);
      LSHR_u32_u32_59_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_73_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_36, konst_72_wire_constant, tmp_var);
      LSHR_u32_u32_73_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_87_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_36, konst_86_wire_constant, tmp_var);
      LSHR_u32_u32_87_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_90_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_36, konst_89_wire_constant, tmp_var);
      LSHR_u32_u32_90_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_217_inst
    process(fetch_val1_129, my_num1_213) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val1_129, my_num1_213, tmp_var);
      LSHR_u64_u64_217_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_240_inst
    process(n_address1_236) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address1_236, konst_239_wire_constant, tmp_var);
      LSHR_u64_u64_240_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_243_inst
    process(address1_102) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_102, konst_242_wire_constant, tmp_var);
      LSHR_u64_u64_243_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_253_inst
    process(n_address1_236) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address1_236, konst_252_wire_constant, tmp_var);
      LSHR_u64_u64_253_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_289_inst
    process(fetch_val2_133, my_num2_285) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val2_133, my_num2_285, tmp_var);
      LSHR_u64_u64_289_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_312_inst
    process(n_address2_308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address2_308, konst_311_wire_constant, tmp_var);
      LSHR_u64_u64_312_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_315_inst
    process(address2_107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_107, konst_314_wire_constant, tmp_var);
      LSHR_u64_u64_315_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_325_inst
    process(n_address2_308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address2_308, konst_324_wire_constant, tmp_var);
      LSHR_u64_u64_325_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_361_inst
    process(fetch_val3_137, my_num3_357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val3_137, my_num3_357, tmp_var);
      LSHR_u64_u64_361_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_384_inst
    process(n_address3_380) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address3_380, konst_383_wire_constant, tmp_var);
      LSHR_u64_u64_384_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_387_inst
    process(address3_112) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address3_112, konst_386_wire_constant, tmp_var);
      LSHR_u64_u64_387_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_397_inst
    process(n_address3_380) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address3_380, konst_396_wire_constant, tmp_var);
      LSHR_u64_u64_397_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_433_inst
    process(fetch_val4_141, my_num4_429) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val4_141, my_num4_429, tmp_var);
      LSHR_u64_u64_433_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_456_inst
    process(n_address4_452) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address4_452, konst_455_wire_constant, tmp_var);
      LSHR_u64_u64_456_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_459_inst
    process(address4_117) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address4_117, konst_458_wire_constant, tmp_var);
      LSHR_u64_u64_459_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_469_inst
    process(n_address4_452) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address4_452, konst_468_wire_constant, tmp_var);
      LSHR_u64_u64_469_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_34_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_34_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_244_inst
    process(LSHR_u64_u64_240_wire, LSHR_u64_u64_243_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_240_wire, LSHR_u64_u64_243_wire, tmp_var);
      NEQ_u64_u1_244_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_316_inst
    process(LSHR_u64_u64_312_wire, LSHR_u64_u64_315_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_312_wire, LSHR_u64_u64_315_wire, tmp_var);
      NEQ_u64_u1_316_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_388_inst
    process(LSHR_u64_u64_384_wire, LSHR_u64_u64_387_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_384_wire, LSHR_u64_u64_387_wire, tmp_var);
      NEQ_u64_u1_388_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_460_inst
    process(LSHR_u64_u64_456_wire, LSHR_u64_u64_459_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_456_wire, LSHR_u64_u64_459_wire, tmp_var);
      NEQ_u64_u1_460_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_40_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(m_factor_36, konst_39_wire_constant, tmp_var);
      m2_factor_41 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_212_inst
    process(SUB_u64_u64_210_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_210_wire, konst_211_wire_constant, tmp_var);
      my_num1_213 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_284_inst
    process(SUB_u64_u64_282_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_282_wire, konst_283_wire_constant, tmp_var);
      my_num2_285 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_356_inst
    process(SUB_u64_u64_354_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_354_wire, konst_355_wire_constant, tmp_var);
      my_num3_357 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_428_inst
    process(SUB_u64_u64_426_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_426_wire, konst_427_wire_constant, tmp_var);
      my_num4_429 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_210_inst
    process(konst_206_wire_constant, AND_u64_u64_209_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_206_wire_constant, AND_u64_u64_209_wire, tmp_var);
      SUB_u64_u64_210_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_282_inst
    process(konst_278_wire_constant, AND_u64_u64_281_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_278_wire_constant, AND_u64_u64_281_wire, tmp_var);
      SUB_u64_u64_282_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_354_inst
    process(konst_350_wire_constant, AND_u64_u64_353_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_350_wire_constant, AND_u64_u64_353_wire, tmp_var);
      SUB_u64_u64_354_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_426_inst
    process(konst_422_wire_constant, AND_u64_u64_425_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_422_wire_constant, AND_u64_u64_425_wire, tmp_var);
      SUB_u64_u64_426_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_172_inst
    process(row1_145, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row1_145, row_in_buffer, tmp_var);
      send_now1_173 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_177_inst
    process(row2_150, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row2_150, row_in_buffer, tmp_var);
      send_now2_178 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_198_inst
    process(n_row1_186, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row1_186, row_in_buffer, tmp_var);
      continue1_199 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_203_inst
    process(n_row2_194, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row2_194, row_in_buffer, tmp_var);
      continue2_204 <= tmp_var; --
    end process;
    -- shared split operator group (60) : array_obj_ref_254_index_offset 
    ApIntAdd_group_60: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_253_scaled;
      array_obj_ref_254_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_254_index_offset_req_0;
      array_obj_ref_254_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_254_index_offset_req_1;
      array_obj_ref_254_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_60_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_60_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : array_obj_ref_326_index_offset 
    ApIntAdd_group_61: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_325_scaled;
      array_obj_ref_326_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_326_index_offset_req_0;
      array_obj_ref_326_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_326_index_offset_req_1;
      array_obj_ref_326_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_61_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_61_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_61",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : array_obj_ref_398_index_offset 
    ApIntAdd_group_62: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_397_scaled;
      array_obj_ref_398_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_398_index_offset_req_0;
      array_obj_ref_398_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_398_index_offset_req_1;
      array_obj_ref_398_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_62_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_62_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_62",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : array_obj_ref_470_index_offset 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_469_scaled;
      array_obj_ref_470_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_470_index_offset_req_0;
      array_obj_ref_470_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_470_index_offset_req_1;
      array_obj_ref_470_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_63_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_63_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : array_obj_ref_61_index_offset 
    ApIntAdd_group_64: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_60_scaled;
      array_obj_ref_61_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_61_index_offset_req_0;
      array_obj_ref_61_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_61_index_offset_req_1;
      array_obj_ref_61_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_64_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_64_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : array_obj_ref_75_index_offset 
    ApIntAdd_group_65: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_74_scaled;
      array_obj_ref_75_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_75_index_offset_req_0;
      array_obj_ref_75_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_75_index_offset_req_1;
      array_obj_ref_75_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_65_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_65_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : array_obj_ref_93_index_offset 
    ApIntAdd_group_66: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_92_scaled;
      array_obj_ref_93_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_93_index_offset_req_0;
      array_obj_ref_93_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_93_index_offset_req_1;
      array_obj_ref_93_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_66_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_66_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared load operator group (0) : ptr_deref_407_load_0 ptr_deref_479_load_0 ptr_deref_52_load_0 ptr_deref_66_load_0 ptr_deref_80_load_0 ptr_deref_98_load_0 ptr_deref_263_load_0 ptr_deref_335_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(111 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 2, 6 => 2, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(7 downto 0) := (7 => 2, 6 => 2, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => true, 1 => true, 2 => false, 3 => false, 4 => false, 5 => false, 6 => true, 7 => true);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 6, 1 => 6, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 6, 7 => 6);
      -- 
    begin -- 
      reqL_unguarded(7) <= ptr_deref_407_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_479_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_52_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_66_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_80_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_98_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_263_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_335_load_0_req_0;
      ptr_deref_407_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_479_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_52_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_66_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_80_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_98_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_263_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_335_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_407_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_479_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_52_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_66_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_80_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_98_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_263_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_335_load_0_req_1;
      ptr_deref_407_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_479_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_52_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_66_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_80_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_98_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_263_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_335_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn2_314_delayed_7_0_331(0);
      guard_vector(1)  <= fn1_254_delayed_7_0_259(0);
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <= fn4_434_delayed_7_0_475(0);
      guard_vector(7)  <= fn3_374_delayed_7_0_403(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_6: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_6", num_slots => 2) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_7: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_7", num_slots => 2) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_407_word_address_0 & ptr_deref_479_word_address_0 & ptr_deref_52_word_address_0 & ptr_deref_66_word_address_0 & ptr_deref_80_word_address_0 & ptr_deref_98_word_address_0 & ptr_deref_263_word_address_0 & ptr_deref_335_word_address_0;
      ptr_deref_407_data_0 <= data_out(511 downto 448);
      ptr_deref_479_data_0 <= data_out(447 downto 384);
      ptr_deref_52_data_0 <= data_out(383 downto 320);
      ptr_deref_66_data_0 <= data_out(319 downto 256);
      ptr_deref_80_data_0 <= data_out(255 downto 192);
      ptr_deref_98_data_0 <= data_out(191 downto 128);
      ptr_deref_263_data_0 <= data_out(127 downto 64);
      ptr_deref_335_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 8,
        tag_length => 4,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_494_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe1_494_inst_req_0;
      WPIPE_input_pipe1_494_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe1_494_inst_req_1;
      WPIPE_input_pipe1_494_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now1_173(0);
      data_in <= var_val1_219;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_input_pipe2_498_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe2_498_inst_req_0;
      WPIPE_input_pipe2_498_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe2_498_inst_req_1;
      WPIPE_input_pipe2_498_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now1_173(0);
      data_in <= var_val2_291;
      input_pipe2_write_1_gI: SplitGuardInterface generic map(name => "input_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "input_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe2_pipe_write_req(0),
          oack => input_pipe2_pipe_write_ack(0),
          odata => input_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_input_pipe3_502_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe3_502_inst_req_0;
      WPIPE_input_pipe3_502_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe3_502_inst_req_1;
      WPIPE_input_pipe3_502_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now1_173(0);
      data_in <= var_val3_363;
      input_pipe3_write_2_gI: SplitGuardInterface generic map(name => "input_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "input_pipe3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe3_pipe_write_req(0),
          oack => input_pipe3_pipe_write_ack(0),
          odata => input_pipe3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_input_pipe4_506_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe4_506_inst_req_0;
      WPIPE_input_pipe4_506_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe4_506_inst_req_1;
      WPIPE_input_pipe4_506_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now2_178(0);
      data_in <= var_val4_435;
      input_pipe4_write_3_gI: SplitGuardInterface generic map(name => "input_pipe4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe4_write_3: OutputPortRevised -- 
        generic map ( name => "input_pipe4", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe4_pipe_write_req(0),
          oack => input_pipe4_pipe_write_ack(0),
          odata => input_pipe4_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(47 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(63 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_3515_start: Boolean;
  signal convolution3D_CP_3515_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_1184_inst_req_0 : boolean;
  signal type_cast_1188_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1184_inst_ack_1 : boolean;
  signal type_cast_1201_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1753_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1184_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1234_inst_ack_1 : boolean;
  signal type_cast_1905_inst_req_0 : boolean;
  signal type_cast_1213_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1234_inst_ack_0 : boolean;
  signal type_cast_1905_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1209_inst_req_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1197_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1234_inst_req_1 : boolean;
  signal type_cast_1226_inst_req_0 : boolean;
  signal addr_of_1964_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1234_inst_req_0 : boolean;
  signal addr_of_1964_final_reg_ack_0 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1184_inst_ack_0 : boolean;
  signal type_cast_1188_inst_ack_1 : boolean;
  signal type_cast_1188_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1222_inst_ack_0 : boolean;
  signal type_cast_1226_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1247_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1247_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1197_inst_ack_1 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1201_inst_ack_0 : boolean;
  signal type_cast_1226_inst_req_1 : boolean;
  signal type_cast_1213_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1247_inst_req_1 : boolean;
  signal addr_of_1964_final_reg_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1222_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1247_inst_ack_1 : boolean;
  signal type_cast_1213_inst_req_1 : boolean;
  signal type_cast_1201_inst_req_1 : boolean;
  signal type_cast_1226_inst_ack_0 : boolean;
  signal type_cast_1772_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1222_inst_req_1 : boolean;
  signal type_cast_1928_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1222_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1209_inst_ack_1 : boolean;
  signal type_cast_1213_inst_ack_1 : boolean;
  signal type_cast_1188_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1209_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1209_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1297_inst_ack_1 : boolean;
  signal array_obj_ref_1963_index_offset_req_1 : boolean;
  signal if_stmt_1875_branch_ack_1 : boolean;
  signal type_cast_1263_inst_req_1 : boolean;
  signal addr_of_1819_final_reg_ack_1 : boolean;
  signal type_cast_1263_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2535_inst_req_0 : boolean;
  signal addr_of_1819_final_reg_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1272_inst_req_0 : boolean;
  signal type_cast_1251_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1272_inst_ack_0 : boolean;
  signal type_cast_1772_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1272_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1272_inst_ack_1 : boolean;
  signal addr_of_1819_final_reg_ack_0 : boolean;
  signal addr_of_1819_final_reg_req_0 : boolean;
  signal type_cast_1251_inst_req_1 : boolean;
  signal type_cast_1923_inst_req_1 : boolean;
  signal type_cast_1288_inst_req_0 : boolean;
  signal type_cast_1288_inst_ack_0 : boolean;
  signal type_cast_1288_inst_req_1 : boolean;
  signal type_cast_1288_inst_ack_1 : boolean;
  signal type_cast_1251_inst_req_0 : boolean;
  signal type_cast_1833_inst_ack_1 : boolean;
  signal type_cast_1251_inst_ack_0 : boolean;
  signal type_cast_1276_inst_req_0 : boolean;
  signal type_cast_1833_inst_ack_0 : boolean;
  signal type_cast_1276_inst_ack_0 : boolean;
  signal type_cast_1923_inst_ack_1 : boolean;
  signal type_cast_1276_inst_req_1 : boolean;
  signal type_cast_1833_inst_req_0 : boolean;
  signal type_cast_1276_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2535_inst_ack_0 : boolean;
  signal if_stmt_1875_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1197_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1284_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1284_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1284_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1284_inst_ack_1 : boolean;
  signal array_obj_ref_1963_index_offset_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1197_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1259_inst_req_1 : boolean;
  signal type_cast_1833_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1259_inst_ack_1 : boolean;
  signal type_cast_1905_inst_ack_1 : boolean;
  signal addr_of_1964_final_reg_req_1 : boolean;
  signal type_cast_1263_inst_req_0 : boolean;
  signal type_cast_1263_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1259_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1259_inst_ack_0 : boolean;
  signal type_cast_1772_inst_ack_0 : boolean;
  signal type_cast_1201_inst_ack_1 : boolean;
  signal type_cast_1301_inst_req_0 : boolean;
  signal type_cast_1301_inst_ack_0 : boolean;
  signal type_cast_1301_inst_req_1 : boolean;
  signal type_cast_1301_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1309_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1309_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1309_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1309_inst_ack_1 : boolean;
  signal type_cast_1313_inst_req_0 : boolean;
  signal type_cast_1313_inst_ack_0 : boolean;
  signal type_cast_1313_inst_req_1 : boolean;
  signal type_cast_1313_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1322_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1322_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1322_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1322_inst_ack_1 : boolean;
  signal type_cast_1326_inst_req_0 : boolean;
  signal type_cast_1326_inst_ack_0 : boolean;
  signal type_cast_1326_inst_req_1 : boolean;
  signal type_cast_1326_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1334_inst_ack_1 : boolean;
  signal type_cast_1338_inst_req_0 : boolean;
  signal type_cast_1338_inst_ack_0 : boolean;
  signal type_cast_1338_inst_req_1 : boolean;
  signal type_cast_1338_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1347_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1347_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1347_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1347_inst_ack_1 : boolean;
  signal type_cast_1351_inst_req_0 : boolean;
  signal type_cast_1351_inst_ack_0 : boolean;
  signal type_cast_1351_inst_req_1 : boolean;
  signal type_cast_1351_inst_ack_1 : boolean;
  signal type_cast_1896_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1359_inst_req_0 : boolean;
  signal type_cast_1829_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1359_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1359_inst_req_1 : boolean;
  signal type_cast_1829_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1359_inst_ack_1 : boolean;
  signal type_cast_1928_inst_ack_1 : boolean;
  signal type_cast_1928_inst_req_1 : boolean;
  signal type_cast_1363_inst_req_0 : boolean;
  signal type_cast_1363_inst_ack_0 : boolean;
  signal type_cast_1923_inst_ack_0 : boolean;
  signal type_cast_1363_inst_req_1 : boolean;
  signal type_cast_1363_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2363_inst_ack_0 : boolean;
  signal if_stmt_1875_branch_req_0 : boolean;
  signal type_cast_1896_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1372_inst_req_0 : boolean;
  signal type_cast_1829_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1372_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1372_inst_req_1 : boolean;
  signal type_cast_1829_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1372_inst_ack_1 : boolean;
  signal array_obj_ref_1818_index_offset_ack_1 : boolean;
  signal array_obj_ref_1818_index_offset_req_1 : boolean;
  signal array_obj_ref_1818_index_offset_ack_0 : boolean;
  signal type_cast_1923_inst_req_0 : boolean;
  signal type_cast_1376_inst_req_0 : boolean;
  signal type_cast_1376_inst_ack_0 : boolean;
  signal type_cast_1376_inst_req_1 : boolean;
  signal type_cast_1376_inst_ack_1 : boolean;
  signal array_obj_ref_1818_index_offset_req_0 : boolean;
  signal type_cast_1385_inst_req_0 : boolean;
  signal type_cast_1385_inst_ack_0 : boolean;
  signal type_cast_1385_inst_req_1 : boolean;
  signal type_cast_1385_inst_ack_1 : boolean;
  signal type_cast_1757_inst_ack_1 : boolean;
  signal type_cast_1757_inst_req_1 : boolean;
  signal type_cast_1389_inst_req_0 : boolean;
  signal type_cast_1389_inst_ack_0 : boolean;
  signal type_cast_1389_inst_req_1 : boolean;
  signal type_cast_1389_inst_ack_1 : boolean;
  signal type_cast_2431_inst_req_1 : boolean;
  signal type_cast_1837_inst_ack_1 : boolean;
  signal ptr_deref_1822_store_0_ack_1 : boolean;
  signal type_cast_1404_inst_req_0 : boolean;
  signal ptr_deref_1822_store_0_req_1 : boolean;
  signal type_cast_1404_inst_ack_0 : boolean;
  signal type_cast_1914_inst_ack_1 : boolean;
  signal type_cast_1404_inst_req_1 : boolean;
  signal type_cast_1404_inst_ack_1 : boolean;
  signal type_cast_1757_inst_ack_0 : boolean;
  signal type_cast_1837_inst_req_1 : boolean;
  signal type_cast_1757_inst_req_0 : boolean;
  signal array_obj_ref_1963_index_offset_ack_0 : boolean;
  signal type_cast_1905_inst_req_1 : boolean;
  signal type_cast_1914_inst_req_1 : boolean;
  signal if_stmt_1412_branch_req_0 : boolean;
  signal if_stmt_1412_branch_ack_1 : boolean;
  signal if_stmt_1412_branch_ack_0 : boolean;
  signal type_cast_1772_inst_req_1 : boolean;
  signal type_cast_1432_inst_req_0 : boolean;
  signal type_cast_1432_inst_ack_0 : boolean;
  signal type_cast_1914_inst_ack_0 : boolean;
  signal type_cast_1432_inst_req_1 : boolean;
  signal type_cast_1432_inst_ack_1 : boolean;
  signal type_cast_2431_inst_ack_1 : boolean;
  signal type_cast_1896_inst_ack_0 : boolean;
  signal type_cast_1914_inst_req_0 : boolean;
  signal type_cast_1448_inst_req_0 : boolean;
  signal type_cast_1448_inst_ack_0 : boolean;
  signal type_cast_1448_inst_req_1 : boolean;
  signal type_cast_1448_inst_ack_1 : boolean;
  signal type_cast_1837_inst_ack_0 : boolean;
  signal type_cast_1837_inst_req_0 : boolean;
  signal type_cast_1457_inst_req_0 : boolean;
  signal ptr_deref_1822_store_0_ack_0 : boolean;
  signal type_cast_1457_inst_ack_0 : boolean;
  signal type_cast_1457_inst_req_1 : boolean;
  signal ptr_deref_1822_store_0_req_0 : boolean;
  signal type_cast_1457_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1753_inst_ack_1 : boolean;
  signal if_stmt_1779_branch_ack_0 : boolean;
  signal type_cast_1467_inst_req_0 : boolean;
  signal type_cast_1467_inst_ack_0 : boolean;
  signal if_stmt_1704_branch_ack_0 : boolean;
  signal type_cast_1467_inst_req_1 : boolean;
  signal type_cast_1467_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1753_inst_req_1 : boolean;
  signal type_cast_1896_inst_req_0 : boolean;
  signal if_stmt_1779_branch_ack_1 : boolean;
  signal if_stmt_1779_branch_req_0 : boolean;
  signal array_obj_ref_1502_index_offset_req_0 : boolean;
  signal array_obj_ref_1502_index_offset_ack_0 : boolean;
  signal array_obj_ref_1502_index_offset_req_1 : boolean;
  signal array_obj_ref_1502_index_offset_ack_1 : boolean;
  signal array_obj_ref_1963_index_offset_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1753_inst_ack_0 : boolean;
  signal type_cast_1928_inst_ack_0 : boolean;
  signal addr_of_1503_final_reg_req_0 : boolean;
  signal addr_of_1503_final_reg_ack_0 : boolean;
  signal addr_of_1503_final_reg_req_1 : boolean;
  signal addr_of_1503_final_reg_ack_1 : boolean;
  signal type_cast_2418_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1506_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1506_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1506_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1506_inst_ack_1 : boolean;
  signal type_cast_1510_inst_req_0 : boolean;
  signal type_cast_1510_inst_ack_0 : boolean;
  signal type_cast_1510_inst_req_1 : boolean;
  signal type_cast_1510_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1519_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1519_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_2308_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1519_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1519_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2363_inst_req_1 : boolean;
  signal type_cast_2533_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_2363_inst_ack_1 : boolean;
  signal type_cast_1523_inst_req_0 : boolean;
  signal type_cast_1523_inst_ack_0 : boolean;
  signal type_cast_1523_inst_req_1 : boolean;
  signal type_cast_1523_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2308_inst_ack_0 : boolean;
  signal type_cast_2483_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1537_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1537_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1537_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1537_inst_ack_1 : boolean;
  signal type_cast_2483_inst_ack_0 : boolean;
  signal type_cast_1541_inst_req_0 : boolean;
  signal type_cast_1541_inst_ack_0 : boolean;
  signal type_cast_1541_inst_req_1 : boolean;
  signal type_cast_1541_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1555_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1555_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_2308_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1555_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1555_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2308_inst_ack_1 : boolean;
  signal type_cast_1559_inst_req_0 : boolean;
  signal type_cast_1559_inst_ack_0 : boolean;
  signal call_stmt_2307_call_req_0 : boolean;
  signal type_cast_1559_inst_req_1 : boolean;
  signal type_cast_1559_inst_ack_1 : boolean;
  signal type_cast_2523_inst_req_1 : boolean;
  signal call_stmt_2307_call_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1573_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1573_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1573_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1573_inst_ack_1 : boolean;
  signal call_stmt_2459_call_req_0 : boolean;
  signal type_cast_1577_inst_req_0 : boolean;
  signal type_cast_1577_inst_ack_0 : boolean;
  signal type_cast_1577_inst_req_1 : boolean;
  signal type_cast_1577_inst_ack_1 : boolean;
  signal type_cast_2427_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_2366_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1591_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1591_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1591_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1591_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2366_inst_ack_0 : boolean;
  signal type_cast_1595_inst_req_0 : boolean;
  signal type_cast_1595_inst_ack_0 : boolean;
  signal type_cast_1595_inst_req_1 : boolean;
  signal type_cast_1595_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2311_inst_req_0 : boolean;
  signal type_cast_2523_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1609_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1609_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1609_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1609_inst_ack_1 : boolean;
  signal type_cast_1613_inst_req_0 : boolean;
  signal type_cast_1613_inst_ack_0 : boolean;
  signal type_cast_1613_inst_req_1 : boolean;
  signal type_cast_1613_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1627_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1627_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1627_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1627_inst_ack_1 : boolean;
  signal type_cast_1631_inst_req_0 : boolean;
  signal type_cast_1631_inst_ack_0 : boolean;
  signal type_cast_1631_inst_req_1 : boolean;
  signal type_cast_1631_inst_ack_1 : boolean;
  signal ptr_deref_1639_store_0_req_0 : boolean;
  signal ptr_deref_1639_store_0_ack_0 : boolean;
  signal ptr_deref_1639_store_0_req_1 : boolean;
  signal ptr_deref_1639_store_0_ack_1 : boolean;
  signal if_stmt_1653_branch_req_0 : boolean;
  signal if_stmt_1653_branch_ack_1 : boolean;
  signal if_stmt_1653_branch_ack_0 : boolean;
  signal if_stmt_1704_branch_req_0 : boolean;
  signal if_stmt_1704_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1967_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1967_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1967_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1967_inst_ack_1 : boolean;
  signal type_cast_1971_inst_req_0 : boolean;
  signal type_cast_1971_inst_ack_0 : boolean;
  signal type_cast_1971_inst_req_1 : boolean;
  signal type_cast_1971_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1980_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1980_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1980_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1980_inst_ack_1 : boolean;
  signal type_cast_1984_inst_req_0 : boolean;
  signal type_cast_1984_inst_ack_0 : boolean;
  signal type_cast_1984_inst_req_1 : boolean;
  signal type_cast_1984_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1998_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1998_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1998_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1998_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_2406_inst_ack_1 : boolean;
  signal type_cast_2002_inst_req_0 : boolean;
  signal type_cast_2002_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2406_inst_req_1 : boolean;
  signal type_cast_2002_inst_req_1 : boolean;
  signal type_cast_2002_inst_ack_1 : boolean;
  signal ptr_deref_2301_store_0_ack_1 : boolean;
  signal ptr_deref_2301_store_0_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2016_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2016_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2016_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2016_inst_ack_1 : boolean;
  signal type_cast_2503_inst_ack_1 : boolean;
  signal type_cast_2503_inst_req_1 : boolean;
  signal type_cast_2418_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_2363_inst_req_0 : boolean;
  signal type_cast_2020_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_2406_inst_ack_0 : boolean;
  signal type_cast_2020_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2406_inst_req_0 : boolean;
  signal type_cast_2020_inst_req_1 : boolean;
  signal type_cast_2020_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2034_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2034_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2034_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2034_inst_ack_1 : boolean;
  signal type_cast_2503_inst_ack_0 : boolean;
  signal type_cast_2503_inst_req_0 : boolean;
  signal type_cast_2418_inst_ack_0 : boolean;
  signal type_cast_2038_inst_req_0 : boolean;
  signal type_cast_2038_inst_ack_0 : boolean;
  signal type_cast_2038_inst_req_1 : boolean;
  signal type_cast_2038_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2538_inst_ack_1 : boolean;
  signal type_cast_2523_inst_ack_0 : boolean;
  signal type_cast_2418_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2052_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2052_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2052_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2052_inst_ack_1 : boolean;
  signal type_cast_2473_inst_ack_1 : boolean;
  signal type_cast_2056_inst_req_0 : boolean;
  signal type_cast_2403_inst_ack_1 : boolean;
  signal type_cast_2056_inst_ack_0 : boolean;
  signal type_cast_2473_inst_req_1 : boolean;
  signal type_cast_2056_inst_req_1 : boolean;
  signal type_cast_2403_inst_req_1 : boolean;
  signal type_cast_2056_inst_ack_1 : boolean;
  signal type_cast_2523_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2538_inst_req_1 : boolean;
  signal type_cast_2341_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2070_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2070_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2070_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2070_inst_ack_1 : boolean;
  signal type_cast_2431_inst_ack_0 : boolean;
  signal type_cast_2533_inst_ack_0 : boolean;
  signal type_cast_2493_inst_ack_1 : boolean;
  signal type_cast_2493_inst_req_1 : boolean;
  signal type_cast_2341_inst_req_1 : boolean;
  signal type_cast_2074_inst_req_0 : boolean;
  signal type_cast_2074_inst_ack_0 : boolean;
  signal type_cast_2074_inst_req_1 : boolean;
  signal type_cast_2403_inst_ack_0 : boolean;
  signal type_cast_2074_inst_ack_1 : boolean;
  signal type_cast_2431_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2088_inst_req_0 : boolean;
  signal type_cast_2403_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2088_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2088_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2088_inst_ack_1 : boolean;
  signal type_cast_2533_inst_req_0 : boolean;
  signal type_cast_2493_inst_ack_0 : boolean;
  signal call_stmt_2414_call_ack_1 : boolean;
  signal call_stmt_2414_call_req_1 : boolean;
  signal type_cast_2341_inst_ack_0 : boolean;
  signal type_cast_2473_inst_ack_0 : boolean;
  signal type_cast_2092_inst_req_0 : boolean;
  signal type_cast_2092_inst_ack_0 : boolean;
  signal type_cast_2473_inst_req_0 : boolean;
  signal type_cast_2092_inst_req_1 : boolean;
  signal type_cast_2092_inst_ack_1 : boolean;
  signal call_stmt_2414_call_ack_0 : boolean;
  signal call_stmt_2414_call_req_0 : boolean;
  signal type_cast_2341_inst_req_0 : boolean;
  signal ptr_deref_2100_store_0_req_0 : boolean;
  signal ptr_deref_2100_store_0_ack_0 : boolean;
  signal WPIPE_output_pipe_2311_inst_ack_1 : boolean;
  signal ptr_deref_2100_store_0_req_1 : boolean;
  signal ptr_deref_2100_store_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2538_inst_ack_0 : boolean;
  signal type_cast_2513_inst_ack_1 : boolean;
  signal type_cast_2331_inst_ack_1 : boolean;
  signal if_stmt_2114_branch_req_0 : boolean;
  signal type_cast_2331_inst_req_1 : boolean;
  signal ptr_deref_2301_store_0_ack_0 : boolean;
  signal if_stmt_2114_branch_ack_1 : boolean;
  signal ptr_deref_2301_store_0_req_0 : boolean;
  signal if_stmt_2114_branch_ack_0 : boolean;
  signal call_stmt_2377_call_ack_1 : boolean;
  signal call_stmt_2377_call_req_1 : boolean;
  signal type_cast_2493_inst_req_0 : boolean;
  signal if_stmt_2165_branch_req_0 : boolean;
  signal call_stmt_2377_call_ack_0 : boolean;
  signal if_stmt_2165_branch_ack_1 : boolean;
  signal call_stmt_2377_call_req_0 : boolean;
  signal if_stmt_2165_branch_ack_0 : boolean;
  signal WPIPE_output_pipe_2311_inst_req_1 : boolean;
  signal call_stmt_2459_call_ack_1 : boolean;
  signal type_cast_2180_inst_req_0 : boolean;
  signal if_stmt_2393_branch_ack_0 : boolean;
  signal type_cast_2180_inst_ack_0 : boolean;
  signal type_cast_2463_inst_ack_1 : boolean;
  signal type_cast_2180_inst_req_1 : boolean;
  signal type_cast_2180_inst_ack_1 : boolean;
  signal type_cast_2513_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2538_inst_req_0 : boolean;
  signal type_cast_2427_inst_ack_1 : boolean;
  signal type_cast_2463_inst_req_1 : boolean;
  signal type_cast_2427_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2218_inst_req_0 : boolean;
  signal if_stmt_2393_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2218_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_2218_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_2218_inst_ack_1 : boolean;
  signal type_cast_2331_inst_ack_0 : boolean;
  signal call_stmt_2459_call_req_1 : boolean;
  signal type_cast_2222_inst_req_0 : boolean;
  signal type_cast_2222_inst_ack_0 : boolean;
  signal type_cast_2222_inst_req_1 : boolean;
  signal if_stmt_2393_branch_req_0 : boolean;
  signal type_cast_2222_inst_ack_1 : boolean;
  signal type_cast_2513_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2410_inst_ack_1 : boolean;
  signal type_cast_2331_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_2410_inst_req_1 : boolean;
  signal type_cast_2463_inst_ack_0 : boolean;
  signal type_cast_2237_inst_req_0 : boolean;
  signal type_cast_2237_inst_ack_0 : boolean;
  signal type_cast_2463_inst_req_0 : boolean;
  signal type_cast_2237_inst_req_1 : boolean;
  signal type_cast_2237_inst_ack_1 : boolean;
  signal type_cast_2533_inst_ack_1 : boolean;
  signal type_cast_2513_inst_req_0 : boolean;
  signal if_stmt_2244_branch_req_0 : boolean;
  signal type_cast_2483_inst_ack_1 : boolean;
  signal if_stmt_2244_branch_ack_1 : boolean;
  signal if_stmt_2244_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2535_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_2366_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_2410_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_2410_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_2366_inst_req_1 : boolean;
  signal type_cast_2427_inst_ack_0 : boolean;
  signal array_obj_ref_2283_index_offset_req_0 : boolean;
  signal array_obj_ref_2283_index_offset_ack_0 : boolean;
  signal call_stmt_2307_call_ack_1 : boolean;
  signal array_obj_ref_2283_index_offset_req_1 : boolean;
  signal array_obj_ref_2283_index_offset_ack_1 : boolean;
  signal call_stmt_2459_call_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2535_inst_req_1 : boolean;
  signal call_stmt_2307_call_req_1 : boolean;
  signal type_cast_2483_inst_req_1 : boolean;
  signal call_stmt_2381_call_ack_1 : boolean;
  signal addr_of_2284_final_reg_req_0 : boolean;
  signal call_stmt_2381_call_req_1 : boolean;
  signal addr_of_2284_final_reg_ack_0 : boolean;
  signal addr_of_2284_final_reg_req_1 : boolean;
  signal addr_of_2284_final_reg_ack_1 : boolean;
  signal WPIPE_output_pipe_2314_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_2314_inst_req_1 : boolean;
  signal WPIPE_output_pipe_2314_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_2314_inst_req_0 : boolean;
  signal call_stmt_2381_call_ack_0 : boolean;
  signal call_stmt_2381_call_req_0 : boolean;
  signal WPIPE_output_pipe_2311_inst_ack_0 : boolean;
  signal ptr_deref_2287_store_0_req_0 : boolean;
  signal ptr_deref_2287_store_0_ack_0 : boolean;
  signal ptr_deref_2287_store_0_req_1 : boolean;
  signal ptr_deref_2287_store_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2541_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2541_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2541_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2541_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2544_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2544_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2544_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2544_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2547_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2547_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2547_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2547_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2550_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2550_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2550_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2550_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2553_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2553_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2553_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2553_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2556_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2556_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2556_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2556_inst_ack_1 : boolean;
  signal phi_stmt_1490_req_1 : boolean;
  signal type_cast_1493_inst_req_0 : boolean;
  signal type_cast_1493_inst_ack_0 : boolean;
  signal type_cast_1493_inst_req_1 : boolean;
  signal type_cast_1493_inst_ack_1 : boolean;
  signal phi_stmt_1490_req_0 : boolean;
  signal phi_stmt_1490_ack_0 : boolean;
  signal phi_stmt_1684_req_1 : boolean;
  signal type_cast_1687_inst_req_0 : boolean;
  signal type_cast_1687_inst_ack_0 : boolean;
  signal type_cast_1687_inst_req_1 : boolean;
  signal type_cast_1687_inst_ack_1 : boolean;
  signal phi_stmt_1684_req_0 : boolean;
  signal phi_stmt_1684_ack_0 : boolean;
  signal phi_stmt_1725_req_0 : boolean;
  signal phi_stmt_1732_req_0 : boolean;
  signal type_cast_1731_inst_req_0 : boolean;
  signal type_cast_1731_inst_ack_0 : boolean;
  signal type_cast_1731_inst_req_1 : boolean;
  signal type_cast_1731_inst_ack_1 : boolean;
  signal phi_stmt_1725_req_1 : boolean;
  signal type_cast_1738_inst_req_0 : boolean;
  signal type_cast_1738_inst_ack_0 : boolean;
  signal type_cast_1738_inst_req_1 : boolean;
  signal type_cast_1738_inst_ack_1 : boolean;
  signal phi_stmt_1732_req_1 : boolean;
  signal phi_stmt_1725_ack_0 : boolean;
  signal phi_stmt_1732_ack_0 : boolean;
  signal type_cast_1789_inst_req_0 : boolean;
  signal type_cast_1789_inst_ack_0 : boolean;
  signal type_cast_1789_inst_req_1 : boolean;
  signal type_cast_1789_inst_ack_1 : boolean;
  signal phi_stmt_1786_req_0 : boolean;
  signal phi_stmt_1786_ack_0 : boolean;
  signal phi_stmt_1951_req_0 : boolean;
  signal type_cast_1957_inst_req_0 : boolean;
  signal type_cast_1957_inst_ack_0 : boolean;
  signal type_cast_1957_inst_req_1 : boolean;
  signal type_cast_1957_inst_ack_1 : boolean;
  signal phi_stmt_1951_req_1 : boolean;
  signal phi_stmt_1951_ack_0 : boolean;
  signal type_cast_2151_inst_req_0 : boolean;
  signal type_cast_2151_inst_ack_0 : boolean;
  signal type_cast_2151_inst_req_1 : boolean;
  signal type_cast_2151_inst_ack_1 : boolean;
  signal phi_stmt_2145_req_1 : boolean;
  signal phi_stmt_2145_req_0 : boolean;
  signal phi_stmt_2145_ack_0 : boolean;
  signal phi_stmt_2197_req_1 : boolean;
  signal phi_stmt_2190_req_1 : boolean;
  signal type_cast_2200_inst_req_0 : boolean;
  signal type_cast_2200_inst_ack_0 : boolean;
  signal type_cast_2200_inst_req_1 : boolean;
  signal type_cast_2200_inst_ack_1 : boolean;
  signal phi_stmt_2197_req_0 : boolean;
  signal type_cast_2193_inst_req_0 : boolean;
  signal type_cast_2193_inst_ack_0 : boolean;
  signal type_cast_2193_inst_req_1 : boolean;
  signal type_cast_2193_inst_ack_1 : boolean;
  signal phi_stmt_2190_req_0 : boolean;
  signal phi_stmt_2190_ack_0 : boolean;
  signal phi_stmt_2197_ack_0 : boolean;
  signal type_cast_2254_inst_req_0 : boolean;
  signal type_cast_2254_inst_ack_0 : boolean;
  signal type_cast_2254_inst_req_1 : boolean;
  signal type_cast_2254_inst_ack_1 : boolean;
  signal phi_stmt_2251_req_0 : boolean;
  signal phi_stmt_2251_ack_0 : boolean;
  signal phi_stmt_2350_req_0 : boolean;
  signal type_cast_2356_inst_req_0 : boolean;
  signal type_cast_2356_inst_ack_0 : boolean;
  signal type_cast_2356_inst_req_1 : boolean;
  signal type_cast_2356_inst_ack_1 : boolean;
  signal phi_stmt_2350_req_1 : boolean;
  signal phi_stmt_2350_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_3515_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_3515_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_3515_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_3515_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_3515: Block -- control-path 
    signal convolution3D_CP_3515_elements: BooleanArray(382 downto 0);
    -- 
  begin -- 
    convolution3D_CP_3515_elements(0) <= convolution3D_CP_3515_start;
    convolution3D_CP_3515_symbol <= convolution3D_CP_3515_elements(313);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411__entry__
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1181/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/branch_block_stmt_1181__entry__
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_Update/cr
      -- 
    rr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => RPIPE_maxpool_input_pipe_1184_inst_req_0); -- 
    cr_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1188_inst_req_1); -- 
    cr_3768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1238_inst_req_1); -- 
    cr_3740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1226_inst_req_1); -- 
    cr_3712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1213_inst_req_1); -- 
    cr_3684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1201_inst_req_1); -- 
    cr_3824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1263_inst_req_1); -- 
    cr_3796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1251_inst_req_1); -- 
    cr_3880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1288_inst_req_1); -- 
    cr_3852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1276_inst_req_1); -- 
    cr_3908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1301_inst_req_1); -- 
    cr_3936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1313_inst_req_1); -- 
    cr_3964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1326_inst_req_1); -- 
    cr_3992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1338_inst_req_1); -- 
    cr_4020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1351_inst_req_1); -- 
    cr_4048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1363_inst_req_1); -- 
    cr_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1376_inst_req_1); -- 
    cr_4090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1385_inst_req_1); -- 
    cr_4104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1389_inst_req_1); -- 
    cr_4118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(0), ack => type_cast_1404_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_update_start_
      -- 
    ra_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1184_inst_ack_0, ack => convolution3D_CP_3515_elements(1)); -- 
    cr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(1), ack => RPIPE_maxpool_input_pipe_1184_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1184_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_Sample/rr
      -- 
    ca_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1184_inst_ack_1, ack => convolution3D_CP_3515_elements(2)); -- 
    rr_3651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(2), ack => type_cast_1188_inst_req_0); -- 
    rr_3665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(2), ack => RPIPE_maxpool_input_pipe_1197_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_Sample/ra
      -- 
    ra_3652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1188_inst_ack_0, ack => convolution3D_CP_3515_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1188_update_completed_
      -- 
    ca_3657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1188_inst_ack_1, ack => convolution3D_CP_3515_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_Sample/$exit
      -- 
    ra_3666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1197_inst_ack_0, ack => convolution3D_CP_3515_elements(5)); -- 
    cr_3670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(5), ack => RPIPE_maxpool_input_pipe_1197_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1197_Update/$exit
      -- 
    ca_3671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1197_inst_ack_1, ack => convolution3D_CP_3515_elements(6)); -- 
    rr_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(6), ack => RPIPE_maxpool_input_pipe_1209_inst_req_0); -- 
    rr_3679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(6), ack => type_cast_1201_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_sample_completed_
      -- 
    ra_3680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_0, ack => convolution3D_CP_3515_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1201_Update/ca
      -- 
    ca_3685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_1, ack => convolution3D_CP_3515_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_Update/$entry
      -- 
    ra_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1209_inst_ack_0, ack => convolution3D_CP_3515_elements(9)); -- 
    cr_3698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(9), ack => RPIPE_maxpool_input_pipe_1209_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1209_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_Sample/$entry
      -- 
    ca_3699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1209_inst_ack_1, ack => convolution3D_CP_3515_elements(10)); -- 
    rr_3707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(10), ack => type_cast_1213_inst_req_0); -- 
    rr_3721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(10), ack => RPIPE_maxpool_input_pipe_1222_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_Sample/$exit
      -- 
    ra_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1213_inst_ack_0, ack => convolution3D_CP_3515_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1213_Update/ca
      -- 
    ca_3713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1213_inst_ack_1, ack => convolution3D_CP_3515_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_update_start_
      -- 
    ra_3722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1222_inst_ack_0, ack => convolution3D_CP_3515_elements(13)); -- 
    cr_3726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(13), ack => RPIPE_maxpool_input_pipe_1222_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1222_update_completed_
      -- 
    ca_3727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1222_inst_ack_1, ack => convolution3D_CP_3515_elements(14)); -- 
    rr_3749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(14), ack => RPIPE_maxpool_input_pipe_1234_inst_req_0); -- 
    rr_3735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(14), ack => type_cast_1226_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_Sample/$exit
      -- 
    ra_3736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1226_inst_ack_0, ack => convolution3D_CP_3515_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1226_update_completed_
      -- 
    ca_3741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1226_inst_ack_1, ack => convolution3D_CP_3515_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_sample_completed_
      -- 
    ra_3750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1234_inst_ack_0, ack => convolution3D_CP_3515_elements(17)); -- 
    cr_3754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(17), ack => RPIPE_maxpool_input_pipe_1234_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1234_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_sample_start_
      -- 
    ca_3755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1234_inst_ack_1, ack => convolution3D_CP_3515_elements(18)); -- 
    rr_3777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(18), ack => RPIPE_maxpool_input_pipe_1247_inst_req_0); -- 
    rr_3763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(18), ack => type_cast_1238_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_Sample/ra
      -- 
    ra_3764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => convolution3D_CP_3515_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1238_update_completed_
      -- 
    ca_3769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => convolution3D_CP_3515_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_sample_completed_
      -- 
    ra_3778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1247_inst_ack_0, ack => convolution3D_CP_3515_elements(21)); -- 
    cr_3782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(21), ack => RPIPE_maxpool_input_pipe_1247_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1247_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_sample_start_
      -- 
    ca_3783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1247_inst_ack_1, ack => convolution3D_CP_3515_elements(22)); -- 
    rr_3791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(22), ack => type_cast_1251_inst_req_0); -- 
    rr_3805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(22), ack => RPIPE_maxpool_input_pipe_1259_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_sample_completed_
      -- 
    ra_3792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_0, ack => convolution3D_CP_3515_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1251_update_completed_
      -- 
    ca_3797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_1, ack => convolution3D_CP_3515_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_Sample/ra
      -- 
    ra_3806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1259_inst_ack_0, ack => convolution3D_CP_3515_elements(25)); -- 
    cr_3810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(25), ack => RPIPE_maxpool_input_pipe_1259_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1259_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_sample_start_
      -- 
    ca_3811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1259_inst_ack_1, ack => convolution3D_CP_3515_elements(26)); -- 
    rr_3833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(26), ack => RPIPE_maxpool_input_pipe_1272_inst_req_0); -- 
    rr_3819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(26), ack => type_cast_1263_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_sample_completed_
      -- 
    ra_3820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1263_inst_ack_0, ack => convolution3D_CP_3515_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1263_update_completed_
      -- 
    ca_3825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1263_inst_ack_1, ack => convolution3D_CP_3515_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_Update/cr
      -- 
    ra_3834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1272_inst_ack_0, ack => convolution3D_CP_3515_elements(29)); -- 
    cr_3838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(29), ack => RPIPE_maxpool_input_pipe_1272_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1272_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_Sample/rr
      -- 
    ca_3839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1272_inst_ack_1, ack => convolution3D_CP_3515_elements(30)); -- 
    rr_3847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(30), ack => type_cast_1276_inst_req_0); -- 
    rr_3861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(30), ack => RPIPE_maxpool_input_pipe_1284_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_Sample/ra
      -- 
    ra_3848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1276_inst_ack_0, ack => convolution3D_CP_3515_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1276_Update/ca
      -- 
    ca_3853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1276_inst_ack_1, ack => convolution3D_CP_3515_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_update_start_
      -- CP-element group 33: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_Update/cr
      -- 
    ra_3862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1284_inst_ack_0, ack => convolution3D_CP_3515_elements(33)); -- 
    cr_3866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(33), ack => RPIPE_maxpool_input_pipe_1284_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1284_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_sample_start_
      -- 
    ca_3867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1284_inst_ack_1, ack => convolution3D_CP_3515_elements(34)); -- 
    rr_3875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(34), ack => type_cast_1288_inst_req_0); -- 
    rr_3889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(34), ack => RPIPE_maxpool_input_pipe_1297_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_Sample/ra
      -- 
    ra_3876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1288_inst_ack_0, ack => convolution3D_CP_3515_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1288_Update/ca
      -- 
    ca_3881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1288_inst_ack_1, ack => convolution3D_CP_3515_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_Update/cr
      -- 
    ra_3890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1297_inst_ack_0, ack => convolution3D_CP_3515_elements(37)); -- 
    cr_3894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(37), ack => RPIPE_maxpool_input_pipe_1297_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1297_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_Sample/rr
      -- 
    ca_3895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1297_inst_ack_1, ack => convolution3D_CP_3515_elements(38)); -- 
    rr_3903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(38), ack => type_cast_1301_inst_req_0); -- 
    rr_3917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(38), ack => RPIPE_maxpool_input_pipe_1309_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_Sample/ra
      -- 
    ra_3904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1301_inst_ack_0, ack => convolution3D_CP_3515_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1301_Update/ca
      -- 
    ca_3909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1301_inst_ack_1, ack => convolution3D_CP_3515_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_Update/cr
      -- 
    ra_3918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1309_inst_ack_0, ack => convolution3D_CP_3515_elements(41)); -- 
    cr_3922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(41), ack => RPIPE_maxpool_input_pipe_1309_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1309_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_Sample/rr
      -- 
    ca_3923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1309_inst_ack_1, ack => convolution3D_CP_3515_elements(42)); -- 
    rr_3931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(42), ack => type_cast_1313_inst_req_0); -- 
    rr_3945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(42), ack => RPIPE_maxpool_input_pipe_1322_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_Sample/ra
      -- 
    ra_3932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1313_inst_ack_0, ack => convolution3D_CP_3515_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1313_Update/ca
      -- 
    ca_3937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1313_inst_ack_1, ack => convolution3D_CP_3515_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_update_start_
      -- CP-element group 45: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_Update/cr
      -- 
    ra_3946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1322_inst_ack_0, ack => convolution3D_CP_3515_elements(45)); -- 
    cr_3950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(45), ack => RPIPE_maxpool_input_pipe_1322_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1322_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_Sample/rr
      -- 
    ca_3951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1322_inst_ack_1, ack => convolution3D_CP_3515_elements(46)); -- 
    rr_3959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(46), ack => type_cast_1326_inst_req_0); -- 
    rr_3973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(46), ack => RPIPE_maxpool_input_pipe_1334_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_Sample/ra
      -- 
    ra_3960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1326_inst_ack_0, ack => convolution3D_CP_3515_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1326_Update/ca
      -- 
    ca_3965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1326_inst_ack_1, ack => convolution3D_CP_3515_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_Update/cr
      -- 
    ra_3974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1334_inst_ack_0, ack => convolution3D_CP_3515_elements(49)); -- 
    cr_3978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(49), ack => RPIPE_maxpool_input_pipe_1334_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1334_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_Sample/rr
      -- 
    ca_3979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1334_inst_ack_1, ack => convolution3D_CP_3515_elements(50)); -- 
    rr_3987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(50), ack => type_cast_1338_inst_req_0); -- 
    rr_4001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(50), ack => RPIPE_maxpool_input_pipe_1347_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_Sample/ra
      -- 
    ra_3988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_0, ack => convolution3D_CP_3515_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1338_Update/ca
      -- 
    ca_3993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_1, ack => convolution3D_CP_3515_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_Update/cr
      -- 
    ra_4002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1347_inst_ack_0, ack => convolution3D_CP_3515_elements(53)); -- 
    cr_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(53), ack => RPIPE_maxpool_input_pipe_1347_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1347_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_Sample/rr
      -- 
    ca_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1347_inst_ack_1, ack => convolution3D_CP_3515_elements(54)); -- 
    rr_4015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(54), ack => type_cast_1351_inst_req_0); -- 
    rr_4029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(54), ack => RPIPE_maxpool_input_pipe_1359_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_Sample/ra
      -- 
    ra_4016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1351_inst_ack_0, ack => convolution3D_CP_3515_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1351_Update/ca
      -- 
    ca_4021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1351_inst_ack_1, ack => convolution3D_CP_3515_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_update_start_
      -- CP-element group 57: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_Update/cr
      -- 
    ra_4030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1359_inst_ack_0, ack => convolution3D_CP_3515_elements(57)); -- 
    cr_4034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(57), ack => RPIPE_maxpool_input_pipe_1359_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1359_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_Sample/rr
      -- 
    ca_4035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1359_inst_ack_1, ack => convolution3D_CP_3515_elements(58)); -- 
    rr_4043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(58), ack => type_cast_1363_inst_req_0); -- 
    rr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(58), ack => RPIPE_maxpool_input_pipe_1372_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_Sample/ra
      -- 
    ra_4044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1363_inst_ack_0, ack => convolution3D_CP_3515_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1363_Update/ca
      -- 
    ca_4049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1363_inst_ack_1, ack => convolution3D_CP_3515_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_update_start_
      -- CP-element group 61: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_Update/cr
      -- 
    ra_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1372_inst_ack_0, ack => convolution3D_CP_3515_elements(61)); -- 
    cr_4062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(61), ack => RPIPE_maxpool_input_pipe_1372_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/RPIPE_maxpool_input_pipe_1372_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_Sample/rr
      -- 
    ca_4063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1372_inst_ack_1, ack => convolution3D_CP_3515_elements(62)); -- 
    rr_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(62), ack => type_cast_1376_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_Sample/ra
      -- 
    ra_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_0, ack => convolution3D_CP_3515_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1376_Update/ca
      -- 
    ca_4077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_1, ack => convolution3D_CP_3515_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	16 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_Sample/rr
      -- 
    rr_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(65), ack => type_cast_1385_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(12) & convolution3D_CP_3515_elements(16);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_Sample/ra
      -- 
    ra_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1385_inst_ack_0, ack => convolution3D_CP_3515_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1385_Update/ca
      -- 
    ca_4091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1385_inst_ack_1, ack => convolution3D_CP_3515_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	24 
    -- CP-element group 68: 	20 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_Sample/rr
      -- 
    rr_4099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(68), ack => type_cast_1389_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(24) & convolution3D_CP_3515_elements(20);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_Sample/ra
      -- 
    ra_4100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1389_inst_ack_0, ack => convolution3D_CP_3515_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1389_Update/ca
      -- 
    ca_4105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1389_inst_ack_1, ack => convolution3D_CP_3515_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	8 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: 	4 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_Sample/rr
      -- 
    rr_4113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(71), ack => type_cast_1404_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(8) & convolution3D_CP_3515_elements(67) & convolution3D_CP_3515_elements(70) & convolution3D_CP_3515_elements(4);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_Sample/ra
      -- 
    ra_4114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1404_inst_ack_0, ack => convolution3D_CP_3515_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/type_cast_1404_Update/ca
      -- 
    ca_4119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1404_inst_ack_1, ack => convolution3D_CP_3515_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	36 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_1181/if_stmt_1412__entry__
      -- CP-element group 74: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411__exit__
      -- CP-element group 74: 	 branch_block_stmt_1181/assign_stmt_1185_to_assign_stmt_1411/$exit
      -- CP-element group 74: 	 branch_block_stmt_1181/if_stmt_1412_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1181/if_stmt_1412_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1181/if_stmt_1412_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1181/if_stmt_1412_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1181/R_cmp383_1413_place
      -- CP-element group 74: 	 branch_block_stmt_1181/if_stmt_1412_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1181/if_stmt_1412_else_link/$entry
      -- 
    branch_req_4127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(74), ack => if_stmt_1412_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(28) & convolution3D_CP_3515_elements(32) & convolution3D_CP_3515_elements(48) & convolution3D_CP_3515_elements(40) & convolution3D_CP_3515_elements(44) & convolution3D_CP_3515_elements(36) & convolution3D_CP_3515_elements(52) & convolution3D_CP_3515_elements(56) & convolution3D_CP_3515_elements(60) & convolution3D_CP_3515_elements(64) & convolution3D_CP_3515_elements(73);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_1181/merge_stmt_1418__exit__
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487__entry__
      -- CP-element group 75: 	 branch_block_stmt_1181/if_stmt_1412_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1181/if_stmt_1412_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1181/entry_bbx_xnph385
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_1181/entry_bbx_xnph385_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/entry_bbx_xnph385_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1181/merge_stmt_1418_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1181/merge_stmt_1418_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1181/merge_stmt_1418_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1181/merge_stmt_1418_PhiAck/dummy
      -- 
    if_choice_transition_4132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1412_branch_ack_1, ack => convolution3D_CP_3515_elements(75)); -- 
    rr_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(75), ack => type_cast_1432_inst_req_0); -- 
    cr_4154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(75), ack => type_cast_1432_inst_req_1); -- 
    rr_4163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(75), ack => type_cast_1448_inst_req_0); -- 
    cr_4168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(75), ack => type_cast_1448_inst_req_1); -- 
    rr_4177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(75), ack => type_cast_1457_inst_req_0); -- 
    cr_4182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(75), ack => type_cast_1457_inst_req_1); -- 
    cr_4196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(75), ack => type_cast_1467_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	320 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_1181/if_stmt_1412_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1181/if_stmt_1412_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1181/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_1181/entry_forx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1181/entry_forx_xend_PhiReq/phi_stmt_1684/$entry
      -- CP-element group 76: 	 branch_block_stmt_1181/entry_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/$entry
      -- 
    else_choice_transition_4136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1412_branch_ack_0, ack => convolution3D_CP_3515_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_Sample/ra
      -- 
    ra_4150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1432_inst_ack_0, ack => convolution3D_CP_3515_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1432_Update/ca
      -- 
    ca_4155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1432_inst_ack_1, ack => convolution3D_CP_3515_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_Sample/ra
      -- 
    ra_4164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1448_inst_ack_0, ack => convolution3D_CP_3515_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1448_Update/ca
      -- 
    ca_4169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1448_inst_ack_1, ack => convolution3D_CP_3515_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_Sample/ra
      -- 
    ra_4178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1457_inst_ack_0, ack => convolution3D_CP_3515_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1457_Update/ca
      -- 
    ca_4183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1457_inst_ack_1, ack => convolution3D_CP_3515_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_Sample/rr
      -- 
    rr_4191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(83), ack => type_cast_1467_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(80) & convolution3D_CP_3515_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_Sample/ra
      -- 
    ra_4192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_0, ack => convolution3D_CP_3515_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/type_cast_1467_Update/ca
      -- 
    ca_4197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1467_inst_ack_1, ack => convolution3D_CP_3515_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	314 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487__exit__
      -- CP-element group 86: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_1181/assign_stmt_1423_to_assign_stmt_1487/$exit
      -- CP-element group 86: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1490/$entry
      -- CP-element group 86: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(78) & convolution3D_CP_3515_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	319 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_Sample/ack
      -- 
    ack_4226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1502_index_offset_ack_0, ack => convolution3D_CP_3515_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	319 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_request/req
      -- 
    ack_4231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1502_index_offset_ack_1, ack => convolution3D_CP_3515_elements(88)); -- 
    req_4240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(88), ack => addr_of_1503_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_request/ack
      -- 
    ack_4241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1503_final_reg_ack_0, ack => convolution3D_CP_3515_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	319 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_complete/ack
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_word_addrgen/root_register_ack
      -- 
    ack_4246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1503_final_reg_ack_1, ack => convolution3D_CP_3515_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	319 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_Update/cr
      -- 
    ra_4255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1506_inst_ack_0, ack => convolution3D_CP_3515_elements(91)); -- 
    cr_4259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(91), ack => RPIPE_maxpool_input_pipe_1506_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_Sample/rr
      -- 
    ca_4260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1506_inst_ack_1, ack => convolution3D_CP_3515_elements(92)); -- 
    rr_4268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(92), ack => type_cast_1510_inst_req_0); -- 
    rr_4282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(92), ack => RPIPE_maxpool_input_pipe_1519_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_Sample/ra
      -- 
    ra_4269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_0, ack => convolution3D_CP_3515_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	319 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_Update/ca
      -- 
    ca_4274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_1, ack => convolution3D_CP_3515_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_update_start_
      -- CP-element group 95: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_Update/cr
      -- 
    ra_4283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1519_inst_ack_0, ack => convolution3D_CP_3515_elements(95)); -- 
    cr_4287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(95), ack => RPIPE_maxpool_input_pipe_1519_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1519_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_Sample/rr
      -- 
    ca_4288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1519_inst_ack_1, ack => convolution3D_CP_3515_elements(96)); -- 
    rr_4296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(96), ack => type_cast_1523_inst_req_0); -- 
    rr_4310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(96), ack => RPIPE_maxpool_input_pipe_1537_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_Sample/ra
      -- 
    ra_4297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1523_inst_ack_0, ack => convolution3D_CP_3515_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	319 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_Update/ca
      -- 
    ca_4302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1523_inst_ack_1, ack => convolution3D_CP_3515_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_update_start_
      -- CP-element group 99: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_Update/cr
      -- 
    ra_4311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1537_inst_ack_0, ack => convolution3D_CP_3515_elements(99)); -- 
    cr_4315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(99), ack => RPIPE_maxpool_input_pipe_1537_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1537_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_Sample/rr
      -- 
    ca_4316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1537_inst_ack_1, ack => convolution3D_CP_3515_elements(100)); -- 
    rr_4324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(100), ack => type_cast_1541_inst_req_0); -- 
    rr_4338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(100), ack => RPIPE_maxpool_input_pipe_1555_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_Sample/ra
      -- 
    ra_4325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1541_inst_ack_0, ack => convolution3D_CP_3515_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	319 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_Update/ca
      -- 
    ca_4330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1541_inst_ack_1, ack => convolution3D_CP_3515_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_update_start_
      -- CP-element group 103: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_Update/cr
      -- 
    ra_4339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1555_inst_ack_0, ack => convolution3D_CP_3515_elements(103)); -- 
    cr_4343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(103), ack => RPIPE_maxpool_input_pipe_1555_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1555_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_Sample/rr
      -- 
    ca_4344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1555_inst_ack_1, ack => convolution3D_CP_3515_elements(104)); -- 
    rr_4352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(104), ack => type_cast_1559_inst_req_0); -- 
    rr_4366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(104), ack => RPIPE_maxpool_input_pipe_1573_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_Sample/ra
      -- 
    ra_4353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1559_inst_ack_0, ack => convolution3D_CP_3515_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	319 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_Update/ca
      -- 
    ca_4358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1559_inst_ack_1, ack => convolution3D_CP_3515_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_update_start_
      -- CP-element group 107: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_Update/cr
      -- 
    ra_4367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1573_inst_ack_0, ack => convolution3D_CP_3515_elements(107)); -- 
    cr_4371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(107), ack => RPIPE_maxpool_input_pipe_1573_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1573_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_Sample/rr
      -- 
    ca_4372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1573_inst_ack_1, ack => convolution3D_CP_3515_elements(108)); -- 
    rr_4380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(108), ack => type_cast_1577_inst_req_0); -- 
    rr_4394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(108), ack => RPIPE_maxpool_input_pipe_1591_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_Sample/ra
      -- 
    ra_4381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_0, ack => convolution3D_CP_3515_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	319 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_Update/ca
      -- 
    ca_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_1, ack => convolution3D_CP_3515_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_update_start_
      -- CP-element group 111: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_Update/cr
      -- 
    ra_4395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1591_inst_ack_0, ack => convolution3D_CP_3515_elements(111)); -- 
    cr_4399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(111), ack => RPIPE_maxpool_input_pipe_1591_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1591_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_Sample/rr
      -- 
    ca_4400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1591_inst_ack_1, ack => convolution3D_CP_3515_elements(112)); -- 
    rr_4408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(112), ack => type_cast_1595_inst_req_0); -- 
    rr_4422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(112), ack => RPIPE_maxpool_input_pipe_1609_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_Sample/ra
      -- 
    ra_4409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1595_inst_ack_0, ack => convolution3D_CP_3515_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	319 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_Update/ca
      -- 
    ca_4414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1595_inst_ack_1, ack => convolution3D_CP_3515_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_update_start_
      -- CP-element group 115: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_Update/cr
      -- 
    ra_4423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1609_inst_ack_0, ack => convolution3D_CP_3515_elements(115)); -- 
    cr_4427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(115), ack => RPIPE_maxpool_input_pipe_1609_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1609_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_Sample/rr
      -- 
    ca_4428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1609_inst_ack_1, ack => convolution3D_CP_3515_elements(116)); -- 
    rr_4436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(116), ack => type_cast_1613_inst_req_0); -- 
    rr_4450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(116), ack => RPIPE_maxpool_input_pipe_1627_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_Sample/ra
      -- 
    ra_4437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_0, ack => convolution3D_CP_3515_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	319 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_Update/ca
      -- 
    ca_4442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_1, ack => convolution3D_CP_3515_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_update_start_
      -- CP-element group 119: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_Update/cr
      -- 
    ra_4451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1627_inst_ack_0, ack => convolution3D_CP_3515_elements(119)); -- 
    cr_4455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(119), ack => RPIPE_maxpool_input_pipe_1627_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1627_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_Sample/rr
      -- 
    ca_4456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1627_inst_ack_1, ack => convolution3D_CP_3515_elements(120)); -- 
    rr_4464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(120), ack => type_cast_1631_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_Sample/ra
      -- 
    ra_4465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1631_inst_ack_0, ack => convolution3D_CP_3515_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	319 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_Update/ca
      -- 
    ca_4470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1631_inst_ack_1, ack => convolution3D_CP_3515_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	106 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/ptr_deref_1639_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/ptr_deref_1639_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/ptr_deref_1639_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/ptr_deref_1639_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/word_access_start/word_0/rr
      -- 
    rr_4508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(123), ack => ptr_deref_1639_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(90) & convolution3D_CP_3515_elements(98) & convolution3D_CP_3515_elements(102) & convolution3D_CP_3515_elements(94) & convolution3D_CP_3515_elements(106) & convolution3D_CP_3515_elements(110) & convolution3D_CP_3515_elements(114) & convolution3D_CP_3515_elements(118) & convolution3D_CP_3515_elements(122);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Sample/word_access_start/word_0/ra
      -- 
    ra_4509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1639_store_0_ack_0, ack => convolution3D_CP_3515_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	319 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Update/word_access_complete/word_0/ca
      -- 
    ca_4520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1639_store_0_ack_1, ack => convolution3D_CP_3515_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	87 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_1181/if_stmt_1653__entry__
      -- CP-element group 126: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652__exit__
      -- CP-element group 126: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/$exit
      -- CP-element group 126: 	 branch_block_stmt_1181/if_stmt_1653_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_1181/if_stmt_1653_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_1181/if_stmt_1653_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_1181/if_stmt_1653_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_1181/R_exitcond28_1654_place
      -- CP-element group 126: 	 branch_block_stmt_1181/if_stmt_1653_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_1181/if_stmt_1653_else_link/$entry
      -- 
    branch_req_4528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(126), ack => if_stmt_1653_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(87) & convolution3D_CP_3515_elements(125);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	321 
    -- CP-element group 127: 	322 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_1181/merge_stmt_1659__exit__
      -- CP-element group 127: 	 branch_block_stmt_1181/assign_stmt_1666_to_assign_stmt_1681__entry__
      -- CP-element group 127: 	 branch_block_stmt_1181/assign_stmt_1666_to_assign_stmt_1681__exit__
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_1181/if_stmt_1653_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_1181/if_stmt_1653_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_1181/assign_stmt_1666_to_assign_stmt_1681/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/assign_stmt_1666_to_assign_stmt_1681/$exit
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_1181/merge_stmt_1659_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_1181/merge_stmt_1659_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/merge_stmt_1659_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_1181/merge_stmt_1659_PhiAck/dummy
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1653_branch_ack_1, ack => convolution3D_CP_3515_elements(127)); -- 
    rr_6079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(127), ack => type_cast_1687_inst_req_0); -- 
    cr_6084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(127), ack => type_cast_1687_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	315 
    -- CP-element group 128: 	316 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_1181/if_stmt_1653_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_1181/if_stmt_1653_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/$entry
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/$entry
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1653_branch_ack_0, ack => convolution3D_CP_3515_elements(128)); -- 
    rr_6025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(128), ack => type_cast_1493_inst_req_0); -- 
    cr_6030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(128), ack => type_cast_1493_inst_req_1); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	325 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	344 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_1181/forx_xend_ifx_xend
      -- CP-element group 129: 	 branch_block_stmt_1181/if_stmt_1704_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_1181/if_stmt_1704_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_1181/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_1181/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_4558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1704_branch_ack_1, ack => convolution3D_CP_3515_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	325 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	326 
    -- CP-element group 130: 	327 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_1181/merge_stmt_1710__exit__
      -- CP-element group 130: 	 branch_block_stmt_1181/assign_stmt_1716_to_assign_stmt_1722__entry__
      -- CP-element group 130: 	 branch_block_stmt_1181/assign_stmt_1716_to_assign_stmt_1722__exit__
      -- CP-element group 130: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_1181/assign_stmt_1716_to_assign_stmt_1722/$exit
      -- CP-element group 130: 	 branch_block_stmt_1181/assign_stmt_1716_to_assign_stmt_1722/$entry
      -- CP-element group 130: 	 branch_block_stmt_1181/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_1181/if_stmt_1704_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_1181/if_stmt_1704_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_1181/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_1181/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_1181/merge_stmt_1710_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_1181/merge_stmt_1710_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_1181/merge_stmt_1710_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_1181/merge_stmt_1710_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/$entry
      -- CP-element group 130: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/$entry
      -- CP-element group 130: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/$entry
      -- 
    else_choice_transition_4562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1704_branch_ack_0, ack => convolution3D_CP_3515_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	339 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_update_start_
      -- 
    ra_4579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1753_inst_ack_0, ack => convolution3D_CP_3515_elements(131)); -- 
    cr_4583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(131), ack => RPIPE_maxpool_input_pipe_1753_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_Update/$exit
      -- 
    ca_4584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1753_inst_ack_1, ack => convolution3D_CP_3515_elements(132)); -- 
    rr_4592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(132), ack => type_cast_1757_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_sample_completed_
      -- 
    ra_4593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1757_inst_ack_0, ack => convolution3D_CP_3515_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	339 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_update_completed_
      -- 
    ca_4598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1757_inst_ack_1, ack => convolution3D_CP_3515_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	339 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_sample_completed_
      -- 
    ra_4607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_0, ack => convolution3D_CP_3515_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	339 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_update_completed_
      -- 
    ca_4612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_1, ack => convolution3D_CP_3515_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_1181/if_stmt_1779__entry__
      -- CP-element group 137: 	 branch_block_stmt_1181/if_stmt_1779_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778__exit__
      -- CP-element group 137: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/$exit
      -- CP-element group 137: 	 branch_block_stmt_1181/R_cmpx_xi_1780_place
      -- CP-element group 137: 	 branch_block_stmt_1181/if_stmt_1779_else_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_1181/if_stmt_1779_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_1181/if_stmt_1779_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_1181/if_stmt_1779_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_1181/if_stmt_1779_eval_test/$entry
      -- 
    branch_req_4620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(137), ack => if_stmt_1779_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(134) & convolution3D_CP_3515_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	329 
    -- CP-element group 138: 	330 
    -- CP-element group 138: 	332 
    -- CP-element group 138: 	333 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_1181/if_stmt_1779_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_1181/if_stmt_1779_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1779_branch_ack_1, ack => convolution3D_CP_3515_elements(138)); -- 
    rr_6141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(138), ack => type_cast_1731_inst_req_0); -- 
    cr_6146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(138), ack => type_cast_1731_inst_req_1); -- 
    rr_6164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(138), ack => type_cast_1738_inst_req_0); -- 
    cr_6169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(138), ack => type_cast_1738_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	340 
    -- CP-element group 139: 	341 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_1181/if_stmt_1779_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_1181/if_stmt_1779_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/$entry
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/$entry
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1779_branch_ack_0, ack => convolution3D_CP_3515_elements(139)); -- 
    rr_6200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(139), ack => type_cast_1789_inst_req_0); -- 
    cr_6205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(139), ack => type_cast_1789_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	343 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_Sample/ack
      -- CP-element group 140: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_sample_complete
      -- 
    ack_4660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1818_index_offset_ack_0, ack => convolution3D_CP_3515_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	343 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_request/req
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_sample_start_
      -- 
    ack_4665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1818_index_offset_ack_1, ack => convolution3D_CP_3515_elements(141)); -- 
    req_4674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(141), ack => addr_of_1819_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_request/ack
      -- CP-element group 142: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_request/$exit
      -- CP-element group 142: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_sample_completed_
      -- 
    ack_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1819_final_reg_ack_0, ack => convolution3D_CP_3515_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	343 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_word_addrgen/root_register_ack
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/word_access_start/word_0/rr
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/ptr_deref_1822_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/ptr_deref_1822_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/ptr_deref_1822_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/ptr_deref_1822_Split/$entry
      -- 
    ack_4680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1819_final_reg_ack_1, ack => convolution3D_CP_3515_elements(143)); -- 
    rr_4718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(143), ack => ptr_deref_1822_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/word_access_start/word_0/ra
      -- CP-element group 144: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Sample/word_access_start/$exit
      -- 
    ra_4719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_0_ack_0, ack => convolution3D_CP_3515_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	343 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Update/word_access_complete/word_0/ca
      -- CP-element group 145: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Update/$exit
      -- 
    ca_4730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1822_store_0_ack_1, ack => convolution3D_CP_3515_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	140 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	344 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_1181/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824__exit__
      -- CP-element group 146: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/$exit
      -- CP-element group 146: 	 branch_block_stmt_1181/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_1181/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(140) & convolution3D_CP_3515_elements(145);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	344 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_sample_completed_
      -- 
    ra_4742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1829_inst_ack_0, ack => convolution3D_CP_3515_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	344 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_update_completed_
      -- 
    ca_4747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1829_inst_ack_1, ack => convolution3D_CP_3515_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	344 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_Sample/$exit
      -- 
    ra_4756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1833_inst_ack_0, ack => convolution3D_CP_3515_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	344 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_Update/$exit
      -- 
    ca_4761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1833_inst_ack_1, ack => convolution3D_CP_3515_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	344 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_Sample/$exit
      -- 
    ra_4770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_0, ack => convolution3D_CP_3515_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	344 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_update_completed_
      -- 
    ca_4775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_1, ack => convolution3D_CP_3515_elements(152)); -- 
    -- CP-element group 153:  branch  join  transition  place  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (10) 
      -- CP-element group 153: 	 branch_block_stmt_1181/R_cmp161379_1876_place
      -- CP-element group 153: 	 branch_block_stmt_1181/if_stmt_1875_else_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_1181/if_stmt_1875__entry__
      -- CP-element group 153: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874__exit__
      -- CP-element group 153: 	 branch_block_stmt_1181/if_stmt_1875_if_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_1181/if_stmt_1875_eval_test/branch_req
      -- CP-element group 153: 	 branch_block_stmt_1181/if_stmt_1875_eval_test/$exit
      -- CP-element group 153: 	 branch_block_stmt_1181/if_stmt_1875_eval_test/$entry
      -- CP-element group 153: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/$exit
      -- CP-element group 153: 	 branch_block_stmt_1181/if_stmt_1875_dead_link/$entry
      -- 
    branch_req_4783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(153), ack => if_stmt_1875_branch_req_0); -- 
    convolution3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(152) & convolution3D_CP_3515_elements(148) & convolution3D_CP_3515_elements(150);
      gj_convolution3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	164 
    -- CP-element group 154: 	166 
    -- CP-element group 154: 	157 
    -- CP-element group 154: 	158 
    -- CP-element group 154: 	159 
    -- CP-element group 154: 	160 
    -- CP-element group 154: 	161 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (36) 
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1181/if_stmt_1875_if_link/if_choice_transition
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/ifx_xend_bbx_xnph
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948__entry__
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1181/merge_stmt_1881__exit__
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1181/if_stmt_1875_if_link/$exit
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1181/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 154: 	 branch_block_stmt_1181/merge_stmt_1881_PhiReqMerge
      -- CP-element group 154: 	 branch_block_stmt_1181/merge_stmt_1881_PhiAck/$entry
      -- CP-element group 154: 	 branch_block_stmt_1181/merge_stmt_1881_PhiAck/$exit
      -- CP-element group 154: 	 branch_block_stmt_1181/merge_stmt_1881_PhiAck/dummy
      -- 
    if_choice_transition_4788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1875_branch_ack_1, ack => convolution3D_CP_3515_elements(154)); -- 
    rr_4819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(154), ack => type_cast_1905_inst_req_0); -- 
    cr_4852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(154), ack => type_cast_1923_inst_req_1); -- 
    cr_4866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(154), ack => type_cast_1928_inst_req_1); -- 
    cr_4810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(154), ack => type_cast_1896_inst_req_1); -- 
    cr_4824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(154), ack => type_cast_1905_inst_req_1); -- 
    cr_4838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(154), ack => type_cast_1914_inst_req_1); -- 
    rr_4833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(154), ack => type_cast_1914_inst_req_0); -- 
    rr_4805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(154), ack => type_cast_1896_inst_req_0); -- 
    -- CP-element group 155:  transition  place  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	354 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1181/ifx_xend_forx_xend215
      -- CP-element group 155: 	 branch_block_stmt_1181/if_stmt_1875_else_link/else_choice_transition
      -- CP-element group 155: 	 branch_block_stmt_1181/if_stmt_1875_else_link/$exit
      -- CP-element group 155: 	 branch_block_stmt_1181/ifx_xend_forx_xend215_PhiReq/$entry
      -- CP-element group 155: 	 branch_block_stmt_1181/ifx_xend_forx_xend215_PhiReq/phi_stmt_2145/$entry
      -- CP-element group 155: 	 branch_block_stmt_1181/ifx_xend_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/$entry
      -- 
    else_choice_transition_4792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1875_branch_ack_0, ack => convolution3D_CP_3515_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_Sample/$exit
      -- 
    ra_4806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1896_inst_ack_0, ack => convolution3D_CP_3515_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1896_Update/$exit
      -- 
    ca_4811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1896_inst_ack_1, ack => convolution3D_CP_3515_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	154 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_Sample/$exit
      -- 
    ra_4820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1905_inst_ack_0, ack => convolution3D_CP_3515_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	154 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	162 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1905_Update/$exit
      -- 
    ca_4825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1905_inst_ack_1, ack => convolution3D_CP_3515_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	154 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_Sample/ra
      -- CP-element group 160: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_sample_completed_
      -- 
    ra_4834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1914_inst_ack_0, ack => convolution3D_CP_3515_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	154 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1914_update_completed_
      -- 
    ca_4839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1914_inst_ack_1, ack => convolution3D_CP_3515_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	157 
    -- CP-element group 162: 	159 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_Sample/rr
      -- CP-element group 162: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_sample_start_
      -- 
    rr_4847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(162), ack => type_cast_1923_inst_req_0); -- 
    convolution3D_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(157) & convolution3D_CP_3515_elements(159) & convolution3D_CP_3515_elements(161);
      gj_convolution3D_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_Sample/ra
      -- CP-element group 163: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_sample_completed_
      -- 
    ra_4848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1923_inst_ack_0, ack => convolution3D_CP_3515_elements(163)); -- 
    -- CP-element group 164:  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	154 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_Sample/rr
      -- CP-element group 164: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_Update/ca
      -- CP-element group 164: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1923_update_completed_
      -- 
    ca_4853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1923_inst_ack_1, ack => convolution3D_CP_3515_elements(164)); -- 
    rr_4861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(164), ack => type_cast_1928_inst_req_0); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_Sample/ra
      -- 
    ra_4862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1928_inst_ack_0, ack => convolution3D_CP_3515_elements(165)); -- 
    -- CP-element group 166:  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	154 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	345 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163
      -- CP-element group 166: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948__exit__
      -- CP-element group 166: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/$exit
      -- CP-element group 166: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_1181/assign_stmt_1887_to_assign_stmt_1948/type_cast_1928_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1951/$entry
      -- CP-element group 166: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/$entry
      -- 
    ca_4867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1928_inst_ack_1, ack => convolution3D_CP_3515_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	350 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	206 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_sample_complete
      -- CP-element group 167: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_Sample/ack
      -- 
    ack_4896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1963_index_offset_ack_0, ack => convolution3D_CP_3515_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	350 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (11) 
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_base_plus_offset/$entry
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_request/req
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_request/$entry
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_offset_calculated
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_root_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_Update/ack
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_base_plus_offset/$exit
      -- 
    ack_4901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1963_index_offset_ack_1, ack => convolution3D_CP_3515_elements(168)); -- 
    req_4910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(168), ack => addr_of_1964_final_reg_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_request/ack
      -- CP-element group 169: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_request/$exit
      -- CP-element group 169: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_sample_completed_
      -- 
    ack_4911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1964_final_reg_ack_0, ack => convolution3D_CP_3515_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	350 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	203 
    -- CP-element group 170:  members (19) 
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_complete/ack
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_complete/$exit
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_word_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_address_resized
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_addr_resize/$entry
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_addr_resize/$exit
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_addr_resize/base_resize_req
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_addr_resize/base_resize_ack
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_word_addrgen/$entry
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_word_addrgen/$exit
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_word_addrgen/root_register_req
      -- CP-element group 170: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_word_addrgen/root_register_ack
      -- 
    ack_4916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1964_final_reg_ack_1, ack => convolution3D_CP_3515_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	350 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_update_start_
      -- CP-element group 171: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_Sample/ra
      -- CP-element group 171: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_Update/cr
      -- 
    ra_4925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1967_inst_ack_0, ack => convolution3D_CP_3515_elements(171)); -- 
    cr_4929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(171), ack => RPIPE_maxpool_input_pipe_1967_inst_req_1); -- 
    -- CP-element group 172:  fork  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: 	175 
    -- CP-element group 172:  members (9) 
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_Update/ca
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_Sample/rr
      -- 
    ca_4930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1967_inst_ack_1, ack => convolution3D_CP_3515_elements(172)); -- 
    rr_4952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(172), ack => RPIPE_maxpool_input_pipe_1980_inst_req_0); -- 
    rr_4938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(172), ack => type_cast_1971_inst_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_Sample/ra
      -- 
    ra_4939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1971_inst_ack_0, ack => convolution3D_CP_3515_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	350 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	203 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_Update/ca
      -- 
    ca_4944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1971_inst_ack_1, ack => convolution3D_CP_3515_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	172 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_update_start_
      -- CP-element group 175: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_Update/cr
      -- 
    ra_4953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1980_inst_ack_0, ack => convolution3D_CP_3515_elements(175)); -- 
    cr_4957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(175), ack => RPIPE_maxpool_input_pipe_1980_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	179 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1980_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_Sample/rr
      -- 
    ca_4958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1980_inst_ack_1, ack => convolution3D_CP_3515_elements(176)); -- 
    rr_4966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(176), ack => type_cast_1984_inst_req_0); -- 
    rr_4980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(176), ack => RPIPE_maxpool_input_pipe_1998_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_Sample/ra
      -- 
    ra_4967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1984_inst_ack_0, ack => convolution3D_CP_3515_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	350 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	203 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_Update/ca
      -- 
    ca_4972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1984_inst_ack_1, ack => convolution3D_CP_3515_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_update_start_
      -- CP-element group 179: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_Update/cr
      -- 
    ra_4981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1998_inst_ack_0, ack => convolution3D_CP_3515_elements(179)); -- 
    cr_4985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(179), ack => RPIPE_maxpool_input_pipe_1998_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1998_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_Sample/rr
      -- 
    ca_4986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1998_inst_ack_1, ack => convolution3D_CP_3515_elements(180)); -- 
    rr_4994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(180), ack => type_cast_2002_inst_req_0); -- 
    rr_5008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(180), ack => RPIPE_maxpool_input_pipe_2016_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_Sample/ra
      -- 
    ra_4995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2002_inst_ack_0, ack => convolution3D_CP_3515_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	350 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	203 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_Update/ca
      -- 
    ca_5000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2002_inst_ack_1, ack => convolution3D_CP_3515_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_update_start_
      -- CP-element group 183: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_Update/cr
      -- 
    ra_5009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2016_inst_ack_0, ack => convolution3D_CP_3515_elements(183)); -- 
    cr_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(183), ack => RPIPE_maxpool_input_pipe_2016_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2016_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_Sample/rr
      -- 
    ca_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2016_inst_ack_1, ack => convolution3D_CP_3515_elements(184)); -- 
    rr_5036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(184), ack => RPIPE_maxpool_input_pipe_2034_inst_req_0); -- 
    rr_5022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(184), ack => type_cast_2020_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_Sample/ra
      -- 
    ra_5023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2020_inst_ack_0, ack => convolution3D_CP_3515_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	350 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	203 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_Update/ca
      -- 
    ca_5028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2020_inst_ack_1, ack => convolution3D_CP_3515_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_update_start_
      -- CP-element group 187: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_Update/cr
      -- 
    ra_5037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2034_inst_ack_0, ack => convolution3D_CP_3515_elements(187)); -- 
    cr_5041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(187), ack => RPIPE_maxpool_input_pipe_2034_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	191 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2034_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_Sample/rr
      -- 
    ca_5042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2034_inst_ack_1, ack => convolution3D_CP_3515_elements(188)); -- 
    rr_5050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(188), ack => type_cast_2038_inst_req_0); -- 
    rr_5064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(188), ack => RPIPE_maxpool_input_pipe_2052_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_Sample/ra
      -- 
    ra_5051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_0, ack => convolution3D_CP_3515_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	350 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	203 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_Update/ca
      -- 
    ca_5056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2038_inst_ack_1, ack => convolution3D_CP_3515_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_update_start_
      -- CP-element group 191: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_Update/cr
      -- 
    ra_5065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2052_inst_ack_0, ack => convolution3D_CP_3515_elements(191)); -- 
    cr_5069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(191), ack => RPIPE_maxpool_input_pipe_2052_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2052_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_Sample/rr
      -- 
    ca_5070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2052_inst_ack_1, ack => convolution3D_CP_3515_elements(192)); -- 
    rr_5078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(192), ack => type_cast_2056_inst_req_0); -- 
    rr_5092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(192), ack => RPIPE_maxpool_input_pipe_2070_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_Sample/ra
      -- 
    ra_5079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2056_inst_ack_0, ack => convolution3D_CP_3515_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	350 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	203 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_Update/ca
      -- 
    ca_5084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2056_inst_ack_1, ack => convolution3D_CP_3515_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_update_start_
      -- CP-element group 195: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_Update/cr
      -- 
    ra_5093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2070_inst_ack_0, ack => convolution3D_CP_3515_elements(195)); -- 
    cr_5097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(195), ack => RPIPE_maxpool_input_pipe_2070_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2070_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_Sample/rr
      -- 
    ca_5098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2070_inst_ack_1, ack => convolution3D_CP_3515_elements(196)); -- 
    rr_5120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(196), ack => RPIPE_maxpool_input_pipe_2088_inst_req_0); -- 
    rr_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(196), ack => type_cast_2074_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_Sample/ra
      -- 
    ra_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2074_inst_ack_0, ack => convolution3D_CP_3515_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	350 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	203 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_Update/ca
      -- 
    ca_5112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2074_inst_ack_1, ack => convolution3D_CP_3515_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_update_start_
      -- CP-element group 199: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_Update/cr
      -- 
    ra_5121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2088_inst_ack_0, ack => convolution3D_CP_3515_elements(199)); -- 
    cr_5125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(199), ack => RPIPE_maxpool_input_pipe_2088_inst_req_1); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_2088_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_Sample/rr
      -- 
    ca_5126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2088_inst_ack_1, ack => convolution3D_CP_3515_elements(200)); -- 
    rr_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(200), ack => type_cast_2092_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_Sample/ra
      -- 
    ra_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2092_inst_ack_0, ack => convolution3D_CP_3515_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	350 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_Update/ca
      -- 
    ca_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2092_inst_ack_1, ack => convolution3D_CP_3515_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	198 
    -- CP-element group 203: 	186 
    -- CP-element group 203: 	202 
    -- CP-element group 203: 	194 
    -- CP-element group 203: 	174 
    -- CP-element group 203: 	182 
    -- CP-element group 203: 	190 
    -- CP-element group 203: 	170 
    -- CP-element group 203: 	178 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (9) 
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/ptr_deref_2100_Split/$entry
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/ptr_deref_2100_Split/$exit
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/ptr_deref_2100_Split/split_req
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/ptr_deref_2100_Split/split_ack
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/word_access_start/$entry
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/word_access_start/word_0/$entry
      -- CP-element group 203: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/word_access_start/word_0/rr
      -- 
    rr_5178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(203), ack => ptr_deref_2100_store_0_req_0); -- 
    convolution3D_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(198) & convolution3D_CP_3515_elements(186) & convolution3D_CP_3515_elements(202) & convolution3D_CP_3515_elements(194) & convolution3D_CP_3515_elements(174) & convolution3D_CP_3515_elements(182) & convolution3D_CP_3515_elements(190) & convolution3D_CP_3515_elements(170) & convolution3D_CP_3515_elements(178);
      gj_convolution3D_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/word_access_start/$exit
      -- CP-element group 204: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/word_access_start/word_0/$exit
      -- CP-element group 204: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Sample/word_access_start/word_0/ra
      -- 
    ra_5179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2100_store_0_ack_0, ack => convolution3D_CP_3515_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	350 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Update/word_access_complete/$exit
      -- CP-element group 205: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Update/word_access_complete/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Update/word_access_complete/word_0/ca
      -- 
    ca_5190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2100_store_0_ack_1, ack => convolution3D_CP_3515_elements(205)); -- 
    -- CP-element group 206:  branch  join  transition  place  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: 	167 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (10) 
      -- CP-element group 206: 	 branch_block_stmt_1181/if_stmt_2114__entry__
      -- CP-element group 206: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/$exit
      -- CP-element group 206: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113__exit__
      -- CP-element group 206: 	 branch_block_stmt_1181/if_stmt_2114_dead_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_1181/if_stmt_2114_eval_test/$entry
      -- CP-element group 206: 	 branch_block_stmt_1181/if_stmt_2114_eval_test/$exit
      -- CP-element group 206: 	 branch_block_stmt_1181/if_stmt_2114_eval_test/branch_req
      -- CP-element group 206: 	 branch_block_stmt_1181/R_exitcond_2115_place
      -- CP-element group 206: 	 branch_block_stmt_1181/if_stmt_2114_if_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_1181/if_stmt_2114_else_link/$entry
      -- 
    branch_req_5198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(206), ack => if_stmt_2114_branch_req_0); -- 
    convolution3D_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(205) & convolution3D_CP_3515_elements(167);
      gj_convolution3D_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	351 
    -- CP-element group 207: 	352 
    -- CP-element group 207:  members (24) 
      -- CP-element group 207: 	 branch_block_stmt_1181/assign_stmt_2127_to_assign_stmt_2142__entry__
      -- CP-element group 207: 	 branch_block_stmt_1181/merge_stmt_2120__exit__
      -- CP-element group 207: 	 branch_block_stmt_1181/assign_stmt_2127_to_assign_stmt_2142__exit__
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 207: 	 branch_block_stmt_1181/if_stmt_2114_if_link/$exit
      -- CP-element group 207: 	 branch_block_stmt_1181/if_stmt_2114_if_link/if_choice_transition
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 207: 	 branch_block_stmt_1181/assign_stmt_2127_to_assign_stmt_2142/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/assign_stmt_2127_to_assign_stmt_2142/$exit
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_1181/merge_stmt_2120_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_1181/merge_stmt_2120_PhiAck/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/merge_stmt_2120_PhiAck/$exit
      -- CP-element group 207: 	 branch_block_stmt_1181/merge_stmt_2120_PhiAck/dummy
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2114_branch_ack_1, ack => convolution3D_CP_3515_elements(207)); -- 
    rr_6308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(207), ack => type_cast_2151_inst_req_0); -- 
    cr_6313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(207), ack => type_cast_2151_inst_req_1); -- 
    -- CP-element group 208:  fork  transition  place  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	346 
    -- CP-element group 208: 	347 
    -- CP-element group 208:  members (12) 
      -- CP-element group 208: 	 branch_block_stmt_1181/if_stmt_2114_else_link/$exit
      -- CP-element group 208: 	 branch_block_stmt_1181/if_stmt_2114_else_link/else_choice_transition
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/$entry
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/$entry
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/$entry
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/$entry
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2114_branch_ack_0, ack => convolution3D_CP_3515_elements(208)); -- 
    rr_6265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(208), ack => type_cast_1957_inst_req_0); -- 
    cr_6270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(208), ack => type_cast_1957_inst_req_1); -- 
    -- CP-element group 209:  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	356 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	375 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_1181/if_stmt_2165_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_1181/if_stmt_2165_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_1181/forx_xend215_ifx_xend227
      -- CP-element group 209: 	 branch_block_stmt_1181/forx_xend215_ifx_xend227_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_1181/forx_xend215_ifx_xend227_PhiReq/$exit
      -- 
    if_choice_transition_5228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2165_branch_ack_1, ack => convolution3D_CP_3515_elements(209)); -- 
    -- CP-element group 210:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	356 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (18) 
      -- CP-element group 210: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187__entry__
      -- CP-element group 210: 	 branch_block_stmt_1181/merge_stmt_2171__exit__
      -- CP-element group 210: 	 branch_block_stmt_1181/if_stmt_2165_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_1181/if_stmt_2165_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_1181/forx_xend215_bbx_xnphx_xi356
      -- CP-element group 210: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/$entry
      -- CP-element group 210: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_update_start_
      -- CP-element group 210: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_Update/cr
      -- CP-element group 210: 	 branch_block_stmt_1181/forx_xend215_bbx_xnphx_xi356_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_1181/forx_xend215_bbx_xnphx_xi356_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_1181/merge_stmt_2171_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_1181/merge_stmt_2171_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_1181/merge_stmt_2171_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_1181/merge_stmt_2171_PhiAck/dummy
      -- 
    else_choice_transition_5232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2165_branch_ack_0, ack => convolution3D_CP_3515_elements(210)); -- 
    rr_5245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(210), ack => type_cast_2180_inst_req_0); -- 
    cr_5250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(210), ack => type_cast_2180_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_Sample/ra
      -- 
    ra_5246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_0, ack => convolution3D_CP_3515_elements(211)); -- 
    -- CP-element group 212:  fork  transition  place  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	358 
    -- CP-element group 212: 	357 
    -- CP-element group 212:  members (11) 
      -- CP-element group 212: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187__exit__
      -- CP-element group 212: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365
      -- CP-element group 212: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/$exit
      -- CP-element group 212: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_1181/assign_stmt_2177_to_assign_stmt_2187/type_cast_2180_Update/ca
      -- CP-element group 212: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/$entry
      -- CP-element group 212: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/$entry
      -- CP-element group 212: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$entry
      -- 
    ca_5251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2180_inst_ack_1, ack => convolution3D_CP_3515_elements(212)); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	370 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_update_start_
      -- CP-element group 213: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_Sample/ra
      -- CP-element group 213: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_Update/cr
      -- 
    ra_5263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2218_inst_ack_0, ack => convolution3D_CP_3515_elements(213)); -- 
    cr_5267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(213), ack => RPIPE_maxpool_input_pipe_2218_inst_req_1); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_Update/ca
      -- CP-element group 214: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_Sample/rr
      -- 
    ca_5268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_2218_inst_ack_1, ack => convolution3D_CP_3515_elements(214)); -- 
    rr_5276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(214), ack => type_cast_2222_inst_req_0); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_Sample/ra
      -- 
    ra_5277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2222_inst_ack_0, ack => convolution3D_CP_3515_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	370 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	219 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_Update/ca
      -- 
    ca_5282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2222_inst_ack_1, ack => convolution3D_CP_3515_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	370 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_Sample/ra
      -- 
    ra_5291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2237_inst_ack_0, ack => convolution3D_CP_3515_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	370 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_Update/ca
      -- 
    ca_5296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2237_inst_ack_1, ack => convolution3D_CP_3515_elements(218)); -- 
    -- CP-element group 219:  branch  join  transition  place  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: 	216 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (10) 
      -- CP-element group 219: 	 branch_block_stmt_1181/if_stmt_2244__entry__
      -- CP-element group 219: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243__exit__
      -- CP-element group 219: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/$exit
      -- CP-element group 219: 	 branch_block_stmt_1181/if_stmt_2244_dead_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_1181/if_stmt_2244_eval_test/$entry
      -- CP-element group 219: 	 branch_block_stmt_1181/if_stmt_2244_eval_test/$exit
      -- CP-element group 219: 	 branch_block_stmt_1181/if_stmt_2244_eval_test/branch_req
      -- CP-element group 219: 	 branch_block_stmt_1181/R_cmpx_xi364_2245_place
      -- CP-element group 219: 	 branch_block_stmt_1181/if_stmt_2244_if_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_1181/if_stmt_2244_else_link/$entry
      -- 
    branch_req_5304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(219), ack => if_stmt_2244_branch_req_0); -- 
    convolution3D_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(218) & convolution3D_CP_3515_elements(216);
      gj_convolution3D_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  place  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	360 
    -- CP-element group 220: 	361 
    -- CP-element group 220: 	363 
    -- CP-element group 220: 	364 
    -- CP-element group 220:  members (20) 
      -- CP-element group 220: 	 branch_block_stmt_1181/if_stmt_2244_if_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_1181/if_stmt_2244_if_link/if_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/Update/cr
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2244_branch_ack_1, ack => convolution3D_CP_3515_elements(220)); -- 
    rr_6381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(220), ack => type_cast_2200_inst_req_0); -- 
    cr_6386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(220), ack => type_cast_2200_inst_req_1); -- 
    rr_6404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(220), ack => type_cast_2193_inst_req_0); -- 
    cr_6409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(220), ack => type_cast_2193_inst_req_1); -- 
    -- CP-element group 221:  fork  transition  place  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	371 
    -- CP-element group 221: 	372 
    -- CP-element group 221:  members (12) 
      -- CP-element group 221: 	 branch_block_stmt_1181/if_stmt_2244_else_link/$exit
      -- CP-element group 221: 	 branch_block_stmt_1181/if_stmt_2244_else_link/else_choice_transition
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/$entry
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/$entry
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/$entry
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Sample/rr
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2244_branch_ack_0, ack => convolution3D_CP_3515_elements(221)); -- 
    rr_6440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(221), ack => type_cast_2254_inst_req_0); -- 
    cr_6445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(221), ack => type_cast_2254_inst_req_1); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	374 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_Sample/ack
      -- 
    ack_5344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2283_index_offset_ack_0, ack => convolution3D_CP_3515_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	374 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_request/req
      -- 
    ack_5349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2283_index_offset_ack_1, ack => convolution3D_CP_3515_elements(223)); -- 
    req_5358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(223), ack => addr_of_2284_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_request/ack
      -- 
    ack_5359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2284_final_reg_ack_0, ack => convolution3D_CP_3515_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	374 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/ptr_deref_2287_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/ptr_deref_2287_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/ptr_deref_2287_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/ptr_deref_2287_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/word_access_start/word_0/rr
      -- 
    ack_5364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2284_final_reg_ack_1, ack => convolution3D_CP_3515_elements(225)); -- 
    rr_5402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(225), ack => ptr_deref_2287_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Sample/word_access_start/word_0/ra
      -- 
    ra_5403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2287_store_0_ack_0, ack => convolution3D_CP_3515_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	374 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Update/word_access_complete/word_0/ca
      -- 
    ca_5414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2287_store_0_ack_1, ack => convolution3D_CP_3515_elements(227)); -- 
    -- CP-element group 228:  join  transition  place  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	375 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_1181/getRemainingElementsx_xexit373_ifx_xend227
      -- CP-element group 228: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289__exit__
      -- CP-element group 228: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/$exit
      -- CP-element group 228: 	 branch_block_stmt_1181/getRemainingElementsx_xexit373_ifx_xend227_PhiReq/$entry
      -- CP-element group 228: 	 branch_block_stmt_1181/getRemainingElementsx_xexit373_ifx_xend227_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(222) & convolution3D_CP_3515_elements(227);
      gj_convolution3D_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	376 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (5) 
      -- CP-element group 229: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/word_access_start/word_0/ra
      -- CP-element group 229: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/word_access_start/word_0/$exit
      -- CP-element group 229: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/word_access_start/$exit
      -- CP-element group 229: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_sample_completed_
      -- 
    ra_5456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2301_store_0_ack_0, ack => convolution3D_CP_3515_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	376 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: 	233 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (18) 
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316__entry__
      -- CP-element group 230: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304__exit__
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_Sample/req
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_Sample/crr
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_update_start_
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/$entry
      -- CP-element group 230: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Update/word_access_complete/word_0/ca
      -- CP-element group 230: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Update/word_access_complete/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Update/word_access_complete/$exit
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_Update/ccr
      -- CP-element group 230: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/$exit
      -- CP-element group 230: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_update_completed_
      -- 
    ca_5467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2301_store_0_ack_1, ack => convolution3D_CP_3515_elements(230)); -- 
    req_5492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(230), ack => WPIPE_output_pipe_2308_inst_req_0); -- 
    crr_5478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(230), ack => call_stmt_2307_call_req_0); -- 
    ccr_5483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(230), ack => call_stmt_2307_call_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_Sample/cra
      -- CP-element group 231: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_sample_completed_
      -- 
    cra_5479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2307_call_ack_0, ack => convolution3D_CP_3515_elements(231)); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	239 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/call_stmt_2307_Update/$exit
      -- 
    cca_5484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2307_call_ack_1, ack => convolution3D_CP_3515_elements(232)); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	230 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_Sample/ack
      -- CP-element group 233: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_Update/req
      -- CP-element group 233: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_update_start_
      -- CP-element group 233: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_sample_completed_
      -- 
    ack_5493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2308_inst_ack_0, ack => convolution3D_CP_3515_elements(233)); -- 
    req_5497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(233), ack => WPIPE_output_pipe_2308_inst_req_1); -- 
    -- CP-element group 234:  transition  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_Update/ack
      -- CP-element group 234: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2308_update_completed_
      -- 
    ack_5498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2308_inst_ack_1, ack => convolution3D_CP_3515_elements(234)); -- 
    req_5506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(234), ack => WPIPE_output_pipe_2311_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_update_start_
      -- CP-element group 235: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_Update/req
      -- CP-element group 235: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_Sample/ack
      -- 
    ack_5507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2311_inst_ack_0, ack => convolution3D_CP_3515_elements(235)); -- 
    req_5511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(235), ack => WPIPE_output_pipe_2311_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2311_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_Sample/$entry
      -- 
    ack_5512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2311_inst_ack_1, ack => convolution3D_CP_3515_elements(236)); -- 
    req_5520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(236), ack => WPIPE_output_pipe_2314_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_Update/req
      -- CP-element group 237: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_update_start_
      -- 
    ack_5521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2314_inst_ack_0, ack => convolution3D_CP_3515_elements(237)); -- 
    req_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(237), ack => WPIPE_output_pipe_2314_inst_req_1); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/WPIPE_output_pipe_2314_update_completed_
      -- 
    ack_5526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_2314_inst_ack_1, ack => convolution3D_CP_3515_elements(238)); -- 
    -- CP-element group 239:  join  fork  transition  place  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	232 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	242 
    -- CP-element group 239: 	243 
    -- CP-element group 239: 	240 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (16) 
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347__entry__
      -- CP-element group 239: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316__exit__
      -- CP-element group 239: 	 branch_block_stmt_1181/call_stmt_2307_to_assign_stmt_2316/$exit
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_Update/cr
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_Sample/rr
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_update_start_
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_Update/cr
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_Sample/rr
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_Sample/$entry
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_update_start_
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_sample_start_
      -- CP-element group 239: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/$entry
      -- 
    cr_5556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(239), ack => type_cast_2341_inst_req_1); -- 
    rr_5551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(239), ack => type_cast_2341_inst_req_0); -- 
    cr_5542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(239), ack => type_cast_2331_inst_req_1); -- 
    rr_5537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(239), ack => type_cast_2331_inst_req_0); -- 
    convolution3D_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(232) & convolution3D_CP_3515_elements(238);
      gj_convolution3D_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_Sample/ra
      -- CP-element group 240: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_sample_completed_
      -- 
    ra_5538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_0, ack => convolution3D_CP_3515_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	244 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_Update/ca
      -- CP-element group 241: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2331_update_completed_
      -- 
    ca_5543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2331_inst_ack_1, ack => convolution3D_CP_3515_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	239 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_Sample/ra
      -- CP-element group 242: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_sample_completed_
      -- 
    ra_5552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_0, ack => convolution3D_CP_3515_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	239 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_Update/ca
      -- CP-element group 243: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/type_cast_2341_update_completed_
      -- 
    ca_5557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2341_inst_ack_1, ack => convolution3D_CP_3515_elements(243)); -- 
    -- CP-element group 244:  join  transition  place  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: 	241 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	377 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody
      -- CP-element group 244: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347__exit__
      -- CP-element group 244: 	 branch_block_stmt_1181/assign_stmt_2323_to_assign_stmt_2347/$exit
      -- CP-element group 244: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- CP-element group 244: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2350/$entry
      -- CP-element group 244: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/$entry
      -- 
    convolution3D_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(243) & convolution3D_CP_3515_elements(241);
      gj_convolution3D_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	382 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_Update/req
      -- CP-element group 245: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_update_start_
      -- CP-element group 245: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_sample_completed_
      -- 
    ack_5569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2363_inst_ack_0, ack => convolution3D_CP_3515_elements(245)); -- 
    req_5573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(245), ack => WPIPE_num_out_pipe_2363_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_update_completed_
      -- 
    ack_5574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2363_inst_ack_1, ack => convolution3D_CP_3515_elements(246)); -- 
    req_5582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(246), ack => WPIPE_num_out_pipe_2366_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_update_start_
      -- CP-element group 247: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_Update/req
      -- 
    ack_5583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2366_inst_ack_0, ack => convolution3D_CP_3515_elements(247)); -- 
    req_5587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(247), ack => WPIPE_num_out_pipe_2366_inst_req_1); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	253 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2366_Update/$exit
      -- 
    ack_5588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_2366_inst_ack_1, ack => convolution3D_CP_3515_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	382 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_Sample/cra
      -- CP-element group 249: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_sample_completed_
      -- 
    cra_5597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2377_call_ack_0, ack => convolution3D_CP_3515_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	382 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	253 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_Update/cca
      -- CP-element group 250: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_update_completed_
      -- 
    cca_5602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2377_call_ack_1, ack => convolution3D_CP_3515_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	382 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_Sample/cra
      -- 
    cra_5611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2381_call_ack_0, ack => convolution3D_CP_3515_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	382 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_Update/cca
      -- CP-element group 252: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_Update/$exit
      -- 
    cca_5616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2381_call_ack_1, ack => convolution3D_CP_3515_elements(252)); -- 
    -- CP-element group 253:  branch  join  transition  place  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	248 
    -- CP-element group 253: 	250 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (10) 
      -- CP-element group 253: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392__exit__
      -- CP-element group 253: 	 branch_block_stmt_1181/if_stmt_2393__entry__
      -- CP-element group 253: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/$exit
      -- CP-element group 253: 	 branch_block_stmt_1181/if_stmt_2393_else_link/$entry
      -- CP-element group 253: 	 branch_block_stmt_1181/if_stmt_2393_if_link/$entry
      -- CP-element group 253: 	 branch_block_stmt_1181/if_stmt_2393_eval_test/branch_req
      -- CP-element group 253: 	 branch_block_stmt_1181/R_exitcond5_2394_place
      -- CP-element group 253: 	 branch_block_stmt_1181/if_stmt_2393_eval_test/$exit
      -- CP-element group 253: 	 branch_block_stmt_1181/if_stmt_2393_eval_test/$entry
      -- CP-element group 253: 	 branch_block_stmt_1181/if_stmt_2393_dead_link/$entry
      -- 
    branch_req_5624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(253), ack => if_stmt_2393_branch_req_0); -- 
    convolution3D_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(248) & convolution3D_CP_3515_elements(250) & convolution3D_CP_3515_elements(252);
      gj_convolution3D_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: 	257 
    -- CP-element group 254: 	258 
    -- CP-element group 254:  members (21) 
      -- CP-element group 254: 	 branch_block_stmt_1181/merge_stmt_2399__exit__
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407__entry__
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_Sample/rr
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_Update/cr
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_Sample/rr
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_update_start_
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/$entry
      -- CP-element group 254: 	 branch_block_stmt_1181/whilex_xbody_whilex_xend
      -- CP-element group 254: 	 branch_block_stmt_1181/if_stmt_2393_if_link/if_choice_transition
      -- CP-element group 254: 	 branch_block_stmt_1181/if_stmt_2393_if_link/$exit
      -- CP-element group 254: 	 branch_block_stmt_1181/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 254: 	 branch_block_stmt_1181/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 254: 	 branch_block_stmt_1181/merge_stmt_2399_PhiReqMerge
      -- CP-element group 254: 	 branch_block_stmt_1181/merge_stmt_2399_PhiAck/$entry
      -- CP-element group 254: 	 branch_block_stmt_1181/merge_stmt_2399_PhiAck/$exit
      -- CP-element group 254: 	 branch_block_stmt_1181/merge_stmt_2399_PhiAck/dummy
      -- 
    if_choice_transition_5629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2393_branch_ack_1, ack => convolution3D_CP_3515_elements(254)); -- 
    rr_5660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(254), ack => RPIPE_input_done_pipe_2406_inst_req_0); -- 
    cr_5651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(254), ack => type_cast_2403_inst_req_1); -- 
    rr_5646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(254), ack => type_cast_2403_inst_req_0); -- 
    -- CP-element group 255:  fork  transition  place  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	378 
    -- CP-element group 255: 	379 
    -- CP-element group 255:  members (12) 
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody
      -- CP-element group 255: 	 branch_block_stmt_1181/if_stmt_2393_else_link/else_choice_transition
      -- CP-element group 255: 	 branch_block_stmt_1181/if_stmt_2393_else_link/$exit
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/$entry
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/$entry
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/$entry
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/$entry
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/Sample/rr
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2393_branch_ack_0, ack => convolution3D_CP_3515_elements(255)); -- 
    rr_6493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(255), ack => type_cast_2356_inst_req_0); -- 
    cr_6498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(255), ack => type_cast_2356_inst_req_1); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_Sample/ra
      -- CP-element group 256: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_sample_completed_
      -- 
    ra_5647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2403_inst_ack_0, ack => convolution3D_CP_3515_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	254 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	260 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_Update/ca
      -- CP-element group 257: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/type_cast_2403_update_completed_
      -- 
    ca_5652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2403_inst_ack_1, ack => convolution3D_CP_3515_elements(257)); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	254 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_Update/cr
      -- CP-element group 258: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_Sample/ra
      -- CP-element group 258: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_update_start_
      -- CP-element group 258: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_sample_completed_
      -- 
    ra_5661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2406_inst_ack_0, ack => convolution3D_CP_3515_elements(258)); -- 
    cr_5665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(258), ack => RPIPE_input_done_pipe_2406_inst_req_1); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_Update/ca
      -- CP-element group 259: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/RPIPE_input_done_pipe_2406_update_completed_
      -- 
    ca_5666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2406_inst_ack_1, ack => convolution3D_CP_3515_elements(259)); -- 
    -- CP-element group 260:  join  transition  place  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	257 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (7) 
      -- CP-element group 260: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407__exit__
      -- CP-element group 260: 	 branch_block_stmt_1181/assign_stmt_2411__entry__
      -- CP-element group 260: 	 branch_block_stmt_1181/assign_stmt_2411/$entry
      -- CP-element group 260: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_1181/assign_stmt_2404_to_assign_stmt_2407/$exit
      -- CP-element group 260: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_Sample/$entry
      -- 
    rr_5677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(260), ack => RPIPE_input_done_pipe_2410_inst_req_0); -- 
    convolution3D_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(257) & convolution3D_CP_3515_elements(259);
      gj_convolution3D_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_update_start_
      -- CP-element group 261: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_Sample/ra
      -- CP-element group 261: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_Sample/$exit
      -- 
    ra_5678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2410_inst_ack_0, ack => convolution3D_CP_3515_elements(261)); -- 
    cr_5682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(261), ack => RPIPE_input_done_pipe_2410_inst_req_1); -- 
    -- CP-element group 262:  fork  transition  place  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	270 
    -- CP-element group 262: 	273 
    -- CP-element group 262: 	263 
    -- CP-element group 262: 	264 
    -- CP-element group 262: 	266 
    -- CP-element group 262: 	267 
    -- CP-element group 262: 	268 
    -- CP-element group 262: 	269 
    -- CP-element group 262:  members (31) 
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459__entry__
      -- CP-element group 262: 	 branch_block_stmt_1181/assign_stmt_2411__exit__
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1181/assign_stmt_2411/$exit
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_Sample/rr
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_Update/ccr
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_Sample/crr
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_Update/ccr
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/$entry
      -- CP-element group 262: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_Update/ca
      -- CP-element group 262: 	 branch_block_stmt_1181/assign_stmt_2411/RPIPE_input_done_pipe_2410_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_Update/$entry
      -- 
    ca_5683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_2410_inst_ack_1, ack => convolution3D_CP_3515_elements(262)); -- 
    cr_5741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(262), ack => type_cast_2431_inst_req_1); -- 
    rr_5722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(262), ack => type_cast_2427_inst_req_0); -- 
    cr_5713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(262), ack => type_cast_2418_inst_req_1); -- 
    rr_5736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(262), ack => type_cast_2431_inst_req_0); -- 
    ccr_5699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(262), ack => call_stmt_2414_call_req_1); -- 
    crr_5694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(262), ack => call_stmt_2414_call_req_0); -- 
    cr_5727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(262), ack => type_cast_2427_inst_req_1); -- 
    ccr_5755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(262), ack => call_stmt_2459_call_req_1); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_Sample/cra
      -- CP-element group 263: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_sample_completed_
      -- 
    cra_5695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2414_call_ack_0, ack => convolution3D_CP_3515_elements(263)); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_Sample/rr
      -- CP-element group 264: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_Update/cca
      -- CP-element group 264: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2414_update_completed_
      -- 
    cca_5700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2414_call_ack_1, ack => convolution3D_CP_3515_elements(264)); -- 
    rr_5708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(264), ack => type_cast_2418_inst_req_0); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_Sample/ra
      -- CP-element group 265: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_sample_completed_
      -- 
    ra_5709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2418_inst_ack_0, ack => convolution3D_CP_3515_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	262 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	274 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_Update/ca
      -- CP-element group 266: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2418_update_completed_
      -- 
    ca_5714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2418_inst_ack_1, ack => convolution3D_CP_3515_elements(266)); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	262 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_Sample/ra
      -- 
    ra_5723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2427_inst_ack_0, ack => convolution3D_CP_3515_elements(267)); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	262 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	271 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2427_Update/$exit
      -- 
    ca_5728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2427_inst_ack_1, ack => convolution3D_CP_3515_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	262 
    -- CP-element group 269: successors 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_Sample/ra
      -- CP-element group 269: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_sample_completed_
      -- 
    ra_5737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_0, ack => convolution3D_CP_3515_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	262 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_Update/ca
      -- CP-element group 270: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/type_cast_2431_update_completed_
      -- 
    ca_5742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_1, ack => convolution3D_CP_3515_elements(270)); -- 
    -- CP-element group 271:  join  transition  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: 	268 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_Sample/crr
      -- CP-element group 271: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_Sample/$entry
      -- 
    crr_5750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(271), ack => call_stmt_2459_call_req_0); -- 
    convolution3D_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(270) & convolution3D_CP_3515_elements(268);
      gj_convolution3D_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_Sample/cra
      -- 
    cra_5751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2459_call_ack_0, ack => convolution3D_CP_3515_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	262 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_Update/cca
      -- CP-element group 273: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/call_stmt_2459_Update/$exit
      -- 
    cca_5756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2459_call_ack_1, ack => convolution3D_CP_3515_elements(273)); -- 
    -- CP-element group 274:  join  fork  transition  place  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: 	266 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274: 	276 
    -- CP-element group 274: 	277 
    -- CP-element group 274: 	278 
    -- CP-element group 274: 	279 
    -- CP-element group 274: 	280 
    -- CP-element group 274: 	281 
    -- CP-element group 274: 	282 
    -- CP-element group 274: 	283 
    -- CP-element group 274: 	284 
    -- CP-element group 274: 	285 
    -- CP-element group 274: 	286 
    -- CP-element group 274: 	287 
    -- CP-element group 274: 	288 
    -- CP-element group 274: 	289 
    -- CP-element group 274: 	290 
    -- CP-element group 274:  members (52) 
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558__entry__
      -- CP-element group 274: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459__exit__
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/call_stmt_2414_to_call_stmt_2459/$exit
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_update_start_
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_update_start_
      -- 
    cr_5870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2533_inst_req_1); -- 
    rr_5795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2483_inst_req_0); -- 
    cr_5856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2523_inst_req_1); -- 
    cr_5828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2503_inst_req_1); -- 
    rr_5823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2503_inst_req_0); -- 
    cr_5786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2473_inst_req_1); -- 
    rr_5851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2523_inst_req_0); -- 
    cr_5814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2493_inst_req_1); -- 
    rr_5865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2533_inst_req_0); -- 
    rr_5781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2473_inst_req_0); -- 
    rr_5809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2493_inst_req_0); -- 
    cr_5842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2513_inst_req_1); -- 
    cr_5772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2463_inst_req_1); -- 
    rr_5767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2463_inst_req_0); -- 
    rr_5837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2513_inst_req_0); -- 
    cr_5800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(274), ack => type_cast_2483_inst_req_1); -- 
    convolution3D_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(273) & convolution3D_CP_3515_elements(266);
      gj_convolution3D_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_Sample/ra
      -- CP-element group 275: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_sample_completed_
      -- 
    ra_5768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2463_inst_ack_0, ack => convolution3D_CP_3515_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	311 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_Update/ca
      -- CP-element group 276: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2463_update_completed_
      -- 
    ca_5773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2463_inst_ack_1, ack => convolution3D_CP_3515_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	274 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_Sample/ra
      -- CP-element group 277: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_sample_completed_
      -- 
    ra_5782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2473_inst_ack_0, ack => convolution3D_CP_3515_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	274 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	308 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_Update/ca
      -- CP-element group 278: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2473_update_completed_
      -- 
    ca_5787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2473_inst_ack_1, ack => convolution3D_CP_3515_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	274 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_sample_completed_
      -- 
    ra_5796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2483_inst_ack_0, ack => convolution3D_CP_3515_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	274 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	305 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2483_Update/ca
      -- 
    ca_5801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2483_inst_ack_1, ack => convolution3D_CP_3515_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	274 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_sample_completed_
      -- 
    ra_5810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2493_inst_ack_0, ack => convolution3D_CP_3515_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	274 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	302 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2493_update_completed_
      -- 
    ca_5815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2493_inst_ack_1, ack => convolution3D_CP_3515_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	274 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_Sample/ra
      -- CP-element group 283: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_sample_completed_
      -- 
    ra_5824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2503_inst_ack_0, ack => convolution3D_CP_3515_elements(283)); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	274 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	299 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_Update/ca
      -- CP-element group 284: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2503_update_completed_
      -- 
    ca_5829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2503_inst_ack_1, ack => convolution3D_CP_3515_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	274 
    -- CP-element group 285: successors 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_Sample/ra
      -- CP-element group 285: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_Sample/$exit
      -- 
    ra_5838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2513_inst_ack_0, ack => convolution3D_CP_3515_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	274 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	296 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_Update/ca
      -- CP-element group 286: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2513_update_completed_
      -- 
    ca_5843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2513_inst_ack_1, ack => convolution3D_CP_3515_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	274 
    -- CP-element group 287: successors 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_Sample/ra
      -- CP-element group 287: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_sample_completed_
      -- 
    ra_5852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2523_inst_ack_0, ack => convolution3D_CP_3515_elements(287)); -- 
    -- CP-element group 288:  transition  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	274 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	293 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_Update/ca
      -- CP-element group 288: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2523_update_completed_
      -- 
    ca_5857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2523_inst_ack_1, ack => convolution3D_CP_3515_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	274 
    -- CP-element group 289: successors 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_sample_completed_
      -- CP-element group 289: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_Sample/ra
      -- CP-element group 289: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_Sample/$exit
      -- 
    ra_5866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2533_inst_ack_0, ack => convolution3D_CP_3515_elements(289)); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	274 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_Update/ca
      -- CP-element group 290: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/type_cast_2533_update_completed_
      -- 
    ca_5871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2533_inst_ack_1, ack => convolution3D_CP_3515_elements(290)); -- 
    req_5879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(290), ack => WPIPE_maxpool_output_pipe_2535_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_update_start_
      -- CP-element group 291: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_Update/req
      -- 
    ack_5880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2535_inst_ack_0, ack => convolution3D_CP_3515_elements(291)); -- 
    req_5884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(291), ack => WPIPE_maxpool_output_pipe_2535_inst_req_1); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2535_Update/ack
      -- 
    ack_5885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2535_inst_ack_1, ack => convolution3D_CP_3515_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	288 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_sample_start_
      -- 
    req_5893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(293), ack => WPIPE_maxpool_output_pipe_2538_inst_req_0); -- 
    convolution3D_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(288) & convolution3D_CP_3515_elements(292);
      gj_convolution3D_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_Update/req
      -- CP-element group 294: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_Sample/ack
      -- CP-element group 294: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_update_start_
      -- CP-element group 294: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_sample_completed_
      -- CP-element group 294: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_Sample/$exit
      -- 
    ack_5894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2538_inst_ack_0, ack => convolution3D_CP_3515_elements(294)); -- 
    req_5898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(294), ack => WPIPE_maxpool_output_pipe_2538_inst_req_1); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_Update/ack
      -- CP-element group 295: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2538_update_completed_
      -- 
    ack_5899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2538_inst_ack_1, ack => convolution3D_CP_3515_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	286 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_Sample/req
      -- 
    req_5907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(296), ack => WPIPE_maxpool_output_pipe_2541_inst_req_0); -- 
    convolution3D_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(286) & convolution3D_CP_3515_elements(295);
      gj_convolution3D_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_update_start_
      -- CP-element group 297: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_Update/req
      -- 
    ack_5908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2541_inst_ack_0, ack => convolution3D_CP_3515_elements(297)); -- 
    req_5912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(297), ack => WPIPE_maxpool_output_pipe_2541_inst_req_1); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2541_Update/ack
      -- 
    ack_5913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2541_inst_ack_1, ack => convolution3D_CP_3515_elements(298)); -- 
    -- CP-element group 299:  join  transition  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	284 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_sample_start_
      -- CP-element group 299: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_Sample/req
      -- 
    req_5921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(299), ack => WPIPE_maxpool_output_pipe_2544_inst_req_0); -- 
    convolution3D_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(284) & convolution3D_CP_3515_elements(298);
      gj_convolution3D_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_update_start_
      -- CP-element group 300: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_Sample/ack
      -- CP-element group 300: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_Update/req
      -- 
    ack_5922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2544_inst_ack_0, ack => convolution3D_CP_3515_elements(300)); -- 
    req_5926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(300), ack => WPIPE_maxpool_output_pipe_2544_inst_req_1); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2544_Update/ack
      -- 
    ack_5927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2544_inst_ack_1, ack => convolution3D_CP_3515_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	282 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_Sample/req
      -- 
    req_5935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(302), ack => WPIPE_maxpool_output_pipe_2547_inst_req_0); -- 
    convolution3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(282) & convolution3D_CP_3515_elements(301);
      gj_convolution3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_update_start_
      -- CP-element group 303: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_Update/req
      -- 
    ack_5936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2547_inst_ack_0, ack => convolution3D_CP_3515_elements(303)); -- 
    req_5940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(303), ack => WPIPE_maxpool_output_pipe_2547_inst_req_1); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2547_Update/ack
      -- 
    ack_5941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2547_inst_ack_1, ack => convolution3D_CP_3515_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	280 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_Sample/req
      -- 
    req_5949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(305), ack => WPIPE_maxpool_output_pipe_2550_inst_req_0); -- 
    convolution3D_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(280) & convolution3D_CP_3515_elements(304);
      gj_convolution3D_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_update_start_
      -- CP-element group 306: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_Sample/ack
      -- CP-element group 306: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_Update/req
      -- 
    ack_5950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2550_inst_ack_0, ack => convolution3D_CP_3515_elements(306)); -- 
    req_5954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(306), ack => WPIPE_maxpool_output_pipe_2550_inst_req_1); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_update_completed_
      -- CP-element group 307: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2550_Update/ack
      -- 
    ack_5955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2550_inst_ack_1, ack => convolution3D_CP_3515_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: 	278 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_Sample/req
      -- 
    req_5963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(308), ack => WPIPE_maxpool_output_pipe_2553_inst_req_0); -- 
    convolution3D_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(307) & convolution3D_CP_3515_elements(278);
      gj_convolution3D_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_update_start_
      -- CP-element group 309: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_Update/req
      -- 
    ack_5964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2553_inst_ack_0, ack => convolution3D_CP_3515_elements(309)); -- 
    req_5968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(309), ack => WPIPE_maxpool_output_pipe_2553_inst_req_1); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2553_Update/ack
      -- 
    ack_5969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2553_inst_ack_1, ack => convolution3D_CP_3515_elements(310)); -- 
    -- CP-element group 311:  join  transition  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: 	276 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_sample_start_
      -- CP-element group 311: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_Sample/$entry
      -- CP-element group 311: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_Sample/req
      -- 
    req_5977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(311), ack => WPIPE_maxpool_output_pipe_2556_inst_req_0); -- 
    convolution3D_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(310) & convolution3D_CP_3515_elements(276);
      gj_convolution3D_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_update_start_
      -- CP-element group 312: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_Sample/ack
      -- CP-element group 312: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_Update/req
      -- 
    ack_5978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2556_inst_ack_0, ack => convolution3D_CP_3515_elements(312)); -- 
    req_5982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(312), ack => WPIPE_maxpool_output_pipe_2556_inst_req_1); -- 
    -- CP-element group 313:  transition  place  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (16) 
      -- CP-element group 313: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558__exit__
      -- CP-element group 313: 	 branch_block_stmt_1181/merge_stmt_2560__exit__
      -- CP-element group 313: 	 branch_block_stmt_1181/branch_block_stmt_1181__exit__
      -- CP-element group 313: 	 branch_block_stmt_1181/$exit
      -- CP-element group 313: 	 branch_block_stmt_1181/return__
      -- CP-element group 313: 	 $exit
      -- CP-element group 313: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/$exit
      -- CP-element group 313: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_1181/assign_stmt_2464_to_assign_stmt_2558/WPIPE_maxpool_output_pipe_2556_Update/ack
      -- CP-element group 313: 	 branch_block_stmt_1181/return___PhiReq/$entry
      -- CP-element group 313: 	 branch_block_stmt_1181/return___PhiReq/$exit
      -- CP-element group 313: 	 branch_block_stmt_1181/merge_stmt_2560_PhiReqMerge
      -- CP-element group 313: 	 branch_block_stmt_1181/merge_stmt_2560_PhiAck/$entry
      -- CP-element group 313: 	 branch_block_stmt_1181/merge_stmt_2560_PhiAck/$exit
      -- CP-element group 313: 	 branch_block_stmt_1181/merge_stmt_2560_PhiAck/dummy
      -- 
    ack_5983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2556_inst_ack_1, ack => convolution3D_CP_3515_elements(313)); -- 
    -- CP-element group 314:  transition  output  delay-element  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	86 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	318 
    -- CP-element group 314:  members (5) 
      -- CP-element group 314: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody_PhiReq/$exit
      -- CP-element group 314: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1490/$exit
      -- CP-element group 314: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/$exit
      -- CP-element group 314: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1496_konst_delay_trans
      -- CP-element group 314: 	 branch_block_stmt_1181/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_req
      -- 
    phi_stmt_1490_req_6006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1490_req_6006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(314), ack => phi_stmt_1490_req_1); -- 
    -- Element group convolution3D_CP_3515_elements(314) is a control-delay.
    cp_element_314_delay: control_delay_element  generic map(name => " 314_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(86), ack => convolution3D_CP_3515_elements(314), clk => clk, reset =>reset);
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	128 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/Sample/ra
      -- 
    ra_6026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1493_inst_ack_0, ack => convolution3D_CP_3515_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	128 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/Update/ca
      -- 
    ca_6031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1493_inst_ack_1, ack => convolution3D_CP_3515_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 317: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/$exit
      -- CP-element group 317: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/$exit
      -- CP-element group 317: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/$exit
      -- CP-element group 317: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_sources/type_cast_1493/SplitProtocol/$exit
      -- CP-element group 317: 	 branch_block_stmt_1181/forx_xbody_forx_xbody_PhiReq/phi_stmt_1490/phi_stmt_1490_req
      -- 
    phi_stmt_1490_req_6032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1490_req_6032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(317), ack => phi_stmt_1490_req_0); -- 
    convolution3D_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(315) & convolution3D_CP_3515_elements(316);
      gj_convolution3D_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  merge  transition  place  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	314 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_1181/merge_stmt_1489_PhiReqMerge
      -- CP-element group 318: 	 branch_block_stmt_1181/merge_stmt_1489_PhiAck/$entry
      -- 
    convolution3D_CP_3515_elements(318) <= OrReduce(convolution3D_CP_3515_elements(314) & convolution3D_CP_3515_elements(317));
    -- CP-element group 319:  fork  transition  place  input  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	91 
    -- CP-element group 319: 	87 
    -- CP-element group 319: 	88 
    -- CP-element group 319: 	90 
    -- CP-element group 319: 	98 
    -- CP-element group 319: 	102 
    -- CP-element group 319: 	94 
    -- CP-element group 319: 	106 
    -- CP-element group 319: 	110 
    -- CP-element group 319: 	114 
    -- CP-element group 319: 	118 
    -- CP-element group 319: 	122 
    -- CP-element group 319: 	125 
    -- CP-element group 319:  members (56) 
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652__entry__
      -- CP-element group 319: 	 branch_block_stmt_1181/merge_stmt_1489__exit__
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_resized_1
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_scaled_1
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_computed_1
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_resize_1/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_resize_1/$exit
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_resize_1/index_resize_req
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_resize_1/index_resize_ack
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_scale_1/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_scale_1/$exit
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_scale_1/scale_rename_req
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_index_scale_1/scale_rename_ack
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_update_start
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_Sample/req
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/array_obj_ref_1502_final_index_sum_regn_Update/req
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_complete/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/addr_of_1503_complete/req
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_sample_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/RPIPE_maxpool_input_pipe_1506_Sample/rr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1510_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1523_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1541_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1559_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1577_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1595_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1613_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/type_cast_1631_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_update_start_
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Update/word_access_complete/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Update/word_access_complete/word_0/$entry
      -- CP-element group 319: 	 branch_block_stmt_1181/assign_stmt_1504_to_assign_stmt_1652/ptr_deref_1639_Update/word_access_complete/word_0/cr
      -- CP-element group 319: 	 branch_block_stmt_1181/merge_stmt_1489_PhiAck/$exit
      -- CP-element group 319: 	 branch_block_stmt_1181/merge_stmt_1489_PhiAck/phi_stmt_1490_ack
      -- 
    phi_stmt_1490_ack_6037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1490_ack_0, ack => convolution3D_CP_3515_elements(319)); -- 
    req_4225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => array_obj_ref_1502_index_offset_req_0); -- 
    req_4230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => array_obj_ref_1502_index_offset_req_1); -- 
    req_4245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => addr_of_1503_final_reg_req_1); -- 
    rr_4254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => RPIPE_maxpool_input_pipe_1506_inst_req_0); -- 
    cr_4273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => type_cast_1510_inst_req_1); -- 
    cr_4301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => type_cast_1523_inst_req_1); -- 
    cr_4329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => type_cast_1541_inst_req_1); -- 
    cr_4357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => type_cast_1559_inst_req_1); -- 
    cr_4385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => type_cast_1577_inst_req_1); -- 
    cr_4413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => type_cast_1595_inst_req_1); -- 
    cr_4441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => type_cast_1613_inst_req_1); -- 
    cr_4469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => type_cast_1631_inst_req_1); -- 
    cr_4519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(319), ack => ptr_deref_1639_store_0_req_1); -- 
    -- CP-element group 320:  transition  output  delay-element  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	76 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	324 
    -- CP-element group 320:  members (5) 
      -- CP-element group 320: 	 branch_block_stmt_1181/entry_forx_xend_PhiReq/$exit
      -- CP-element group 320: 	 branch_block_stmt_1181/entry_forx_xend_PhiReq/phi_stmt_1684/$exit
      -- CP-element group 320: 	 branch_block_stmt_1181/entry_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/$exit
      -- CP-element group 320: 	 branch_block_stmt_1181/entry_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1690_konst_delay_trans
      -- CP-element group 320: 	 branch_block_stmt_1181/entry_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_req
      -- 
    phi_stmt_1684_req_6060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1684_req_6060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(320), ack => phi_stmt_1684_req_1); -- 
    -- Element group convolution3D_CP_3515_elements(320) is a control-delay.
    cp_element_320_delay: control_delay_element  generic map(name => " 320_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(76), ack => convolution3D_CP_3515_elements(320), clk => clk, reset =>reset);
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	127 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/Sample/ra
      -- 
    ra_6080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1687_inst_ack_0, ack => convolution3D_CP_3515_elements(321)); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	127 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (2) 
      -- CP-element group 322: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/Update/ca
      -- 
    ca_6085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1687_inst_ack_1, ack => convolution3D_CP_3515_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 323: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/$exit
      -- CP-element group 323: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/$exit
      -- CP-element group 323: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/$exit
      -- CP-element group 323: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_sources/type_cast_1687/SplitProtocol/$exit
      -- CP-element group 323: 	 branch_block_stmt_1181/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1684/phi_stmt_1684_req
      -- 
    phi_stmt_1684_req_6086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1684_req_6086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(323), ack => phi_stmt_1684_req_0); -- 
    convolution3D_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(321) & convolution3D_CP_3515_elements(322);
      gj_convolution3D_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  merge  transition  place  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: 	320 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (2) 
      -- CP-element group 324: 	 branch_block_stmt_1181/merge_stmt_1683_PhiReqMerge
      -- CP-element group 324: 	 branch_block_stmt_1181/merge_stmt_1683_PhiAck/$entry
      -- 
    convolution3D_CP_3515_elements(324) <= OrReduce(convolution3D_CP_3515_elements(323) & convolution3D_CP_3515_elements(320));
    -- CP-element group 325:  branch  transition  place  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	129 
    -- CP-element group 325: 	130 
    -- CP-element group 325:  members (15) 
      -- CP-element group 325: 	 branch_block_stmt_1181/assign_stmt_1697_to_assign_stmt_1703__exit__
      -- CP-element group 325: 	 branch_block_stmt_1181/merge_stmt_1683__exit__
      -- CP-element group 325: 	 branch_block_stmt_1181/if_stmt_1704__entry__
      -- CP-element group 325: 	 branch_block_stmt_1181/assign_stmt_1697_to_assign_stmt_1703__entry__
      -- CP-element group 325: 	 branch_block_stmt_1181/if_stmt_1704_else_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_1181/assign_stmt_1697_to_assign_stmt_1703/$entry
      -- CP-element group 325: 	 branch_block_stmt_1181/assign_stmt_1697_to_assign_stmt_1703/$exit
      -- CP-element group 325: 	 branch_block_stmt_1181/if_stmt_1704_dead_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_1181/if_stmt_1704_eval_test/$entry
      -- CP-element group 325: 	 branch_block_stmt_1181/if_stmt_1704_eval_test/$exit
      -- CP-element group 325: 	 branch_block_stmt_1181/if_stmt_1704_eval_test/branch_req
      -- CP-element group 325: 	 branch_block_stmt_1181/R_tobool_1705_place
      -- CP-element group 325: 	 branch_block_stmt_1181/if_stmt_1704_if_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_1181/merge_stmt_1683_PhiAck/$exit
      -- CP-element group 325: 	 branch_block_stmt_1181/merge_stmt_1683_PhiAck/phi_stmt_1684_ack
      -- 
    phi_stmt_1684_ack_6091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1684_ack_0, ack => convolution3D_CP_3515_elements(325)); -- 
    branch_req_4553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(325), ack => if_stmt_1704_branch_req_0); -- 
    -- CP-element group 326:  transition  output  delay-element  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	130 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (4) 
      -- CP-element group 326: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/$exit
      -- CP-element group 326: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/$exit
      -- CP-element group 326: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1729_konst_delay_trans
      -- CP-element group 326: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_req
      -- 
    phi_stmt_1725_req_6114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1725_req_6114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(326), ack => phi_stmt_1725_req_0); -- 
    -- Element group convolution3D_CP_3515_elements(326) is a control-delay.
    cp_element_326_delay: control_delay_element  generic map(name => " 326_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(130), ack => convolution3D_CP_3515_elements(326), clk => clk, reset =>reset);
    -- CP-element group 327:  transition  output  delay-element  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	130 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (4) 
      -- CP-element group 327: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/$exit
      -- CP-element group 327: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/$exit
      -- CP-element group 327: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1736_konst_delay_trans
      -- CP-element group 327: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_req
      -- 
    phi_stmt_1732_req_6122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1732_req_6122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(327), ack => phi_stmt_1732_req_0); -- 
    -- Element group convolution3D_CP_3515_elements(327) is a control-delay.
    cp_element_327_delay: control_delay_element  generic map(name => " 327_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(130), ack => convolution3D_CP_3515_elements(327), clk => clk, reset =>reset);
    -- CP-element group 328:  join  transition  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	336 
    -- CP-element group 328:  members (1) 
      -- CP-element group 328: 	 branch_block_stmt_1181/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(326) & convolution3D_CP_3515_elements(327);
      gj_convolution3D_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	138 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (2) 
      -- CP-element group 329: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/Sample/ra
      -- 
    ra_6142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_0, ack => convolution3D_CP_3515_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	138 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	331 
    -- CP-element group 330:  members (2) 
      -- CP-element group 330: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/Update/ca
      -- 
    ca_6147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1731_inst_ack_1, ack => convolution3D_CP_3515_elements(330)); -- 
    -- CP-element group 331:  join  transition  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: 	330 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	335 
    -- CP-element group 331:  members (5) 
      -- CP-element group 331: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/$exit
      -- CP-element group 331: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/$exit
      -- CP-element group 331: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/$exit
      -- CP-element group 331: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_sources/type_cast_1731/SplitProtocol/$exit
      -- CP-element group 331: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1725/phi_stmt_1725_req
      -- 
    phi_stmt_1725_req_6148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1725_req_6148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(331), ack => phi_stmt_1725_req_1); -- 
    convolution3D_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(329) & convolution3D_CP_3515_elements(330);
      gj_convolution3D_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	138 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	334 
    -- CP-element group 332:  members (2) 
      -- CP-element group 332: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/Sample/$exit
      -- CP-element group 332: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/Sample/ra
      -- 
    ra_6165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1738_inst_ack_0, ack => convolution3D_CP_3515_elements(332)); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	138 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (2) 
      -- CP-element group 333: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/Update/ca
      -- 
    ca_6170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1738_inst_ack_1, ack => convolution3D_CP_3515_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	332 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (5) 
      -- CP-element group 334: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/$exit
      -- CP-element group 334: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/$exit
      -- CP-element group 334: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/$exit
      -- CP-element group 334: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_sources/type_cast_1738/SplitProtocol/$exit
      -- CP-element group 334: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1732/phi_stmt_1732_req
      -- 
    phi_stmt_1732_req_6171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1732_req_6171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(334), ack => phi_stmt_1732_req_1); -- 
    convolution3D_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(332) & convolution3D_CP_3515_elements(333);
      gj_convolution3D_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	331 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (1) 
      -- CP-element group 335: 	 branch_block_stmt_1181/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(331) & convolution3D_CP_3515_elements(334);
      gj_convolution3D_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  merge  fork  transition  place  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	328 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336: 	338 
    -- CP-element group 336:  members (2) 
      -- CP-element group 336: 	 branch_block_stmt_1181/merge_stmt_1724_PhiReqMerge
      -- CP-element group 336: 	 branch_block_stmt_1181/merge_stmt_1724_PhiAck/$entry
      -- 
    convolution3D_CP_3515_elements(336) <= OrReduce(convolution3D_CP_3515_elements(328) & convolution3D_CP_3515_elements(335));
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	339 
    -- CP-element group 337:  members (1) 
      -- CP-element group 337: 	 branch_block_stmt_1181/merge_stmt_1724_PhiAck/phi_stmt_1725_ack
      -- 
    phi_stmt_1725_ack_6176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1725_ack_0, ack => convolution3D_CP_3515_elements(337)); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (1) 
      -- CP-element group 338: 	 branch_block_stmt_1181/merge_stmt_1724_PhiAck/phi_stmt_1732_ack
      -- 
    phi_stmt_1732_ack_6177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1732_ack_0, ack => convolution3D_CP_3515_elements(338)); -- 
    -- CP-element group 339:  join  fork  transition  place  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	134 
    -- CP-element group 339: 	135 
    -- CP-element group 339: 	136 
    -- CP-element group 339: 	131 
    -- CP-element group 339:  members (16) 
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_Sample/rr
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_1181/merge_stmt_1724__exit__
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778__entry__
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/RPIPE_maxpool_input_pipe_1753_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_Sample/rr
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_update_start_
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_Update/cr
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/$entry
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1772_Update/cr
      -- CP-element group 339: 	 branch_block_stmt_1181/assign_stmt_1745_to_assign_stmt_1778/type_cast_1757_update_start_
      -- CP-element group 339: 	 branch_block_stmt_1181/merge_stmt_1724_PhiAck/$exit
      -- 
    rr_4578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(339), ack => RPIPE_maxpool_input_pipe_1753_inst_req_0); -- 
    rr_4606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(339), ack => type_cast_1772_inst_req_0); -- 
    cr_4597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(339), ack => type_cast_1757_inst_req_1); -- 
    cr_4611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(339), ack => type_cast_1772_inst_req_1); -- 
    convolution3D_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(337) & convolution3D_CP_3515_elements(338);
      gj_convolution3D_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	139 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	342 
    -- CP-element group 340:  members (2) 
      -- CP-element group 340: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/Sample/ra
      -- 
    ra_6201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1789_inst_ack_0, ack => convolution3D_CP_3515_elements(340)); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	139 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (2) 
      -- CP-element group 341: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/Update/ca
      -- 
    ca_6206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1789_inst_ack_1, ack => convolution3D_CP_3515_elements(341)); -- 
    -- CP-element group 342:  join  transition  place  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (8) 
      -- CP-element group 342: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 342: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/$exit
      -- CP-element group 342: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/$exit
      -- CP-element group 342: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/$exit
      -- CP-element group 342: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_sources/type_cast_1789/SplitProtocol/$exit
      -- CP-element group 342: 	 branch_block_stmt_1181/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1786/phi_stmt_1786_req
      -- CP-element group 342: 	 branch_block_stmt_1181/merge_stmt_1785_PhiReqMerge
      -- CP-element group 342: 	 branch_block_stmt_1181/merge_stmt_1785_PhiAck/$entry
      -- 
    phi_stmt_1786_req_6207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1786_req_6207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(342), ack => phi_stmt_1786_req_0); -- 
    convolution3D_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(340) & convolution3D_CP_3515_elements(341);
      gj_convolution3D_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	140 
    -- CP-element group 343: 	141 
    -- CP-element group 343: 	145 
    -- CP-element group 343: 	143 
    -- CP-element group 343:  members (29) 
      -- CP-element group 343: 	 branch_block_stmt_1181/merge_stmt_1785__exit__
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_complete/req
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_complete/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824__entry__
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_update_start_
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_Update/req
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_Sample/req
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_final_index_sum_regn_update_start
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_scale_1/scale_rename_ack
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_scale_1/scale_rename_req
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_scale_1/$exit
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_scale_1/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_resize_1/index_resize_ack
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_resize_1/index_resize_req
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_resize_1/$exit
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_resize_1/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_computed_1
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Update/word_access_complete/word_0/cr
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_scaled_1
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/array_obj_ref_1818_index_resized_1
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Update/word_access_complete/word_0/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Update/word_access_complete/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/ptr_deref_1822_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/addr_of_1819_update_start_
      -- CP-element group 343: 	 branch_block_stmt_1181/assign_stmt_1796_to_assign_stmt_1824/$entry
      -- CP-element group 343: 	 branch_block_stmt_1181/merge_stmt_1785_PhiAck/$exit
      -- CP-element group 343: 	 branch_block_stmt_1181/merge_stmt_1785_PhiAck/phi_stmt_1786_ack
      -- 
    phi_stmt_1786_ack_6212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1786_ack_0, ack => convolution3D_CP_3515_elements(343)); -- 
    req_4679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(343), ack => addr_of_1819_final_reg_req_1); -- 
    req_4664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(343), ack => array_obj_ref_1818_index_offset_req_1); -- 
    req_4659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(343), ack => array_obj_ref_1818_index_offset_req_0); -- 
    cr_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(343), ack => ptr_deref_1822_store_0_req_1); -- 
    -- CP-element group 344:  merge  fork  transition  place  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	146 
    -- CP-element group 344: 	129 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	147 
    -- CP-element group 344: 	151 
    -- CP-element group 344: 	152 
    -- CP-element group 344: 	148 
    -- CP-element group 344: 	149 
    -- CP-element group 344: 	150 
    -- CP-element group 344:  members (25) 
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_update_start_
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_update_start_
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_Sample/rr
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874__entry__
      -- CP-element group 344: 	 branch_block_stmt_1181/merge_stmt_1826__exit__
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1833_Update/cr
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_Update/cr
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_Sample/rr
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_update_start_
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1829_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/$entry
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_Update/cr
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_Sample/rr
      -- CP-element group 344: 	 branch_block_stmt_1181/assign_stmt_1830_to_assign_stmt_1874/type_cast_1837_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_1181/merge_stmt_1826_PhiReqMerge
      -- CP-element group 344: 	 branch_block_stmt_1181/merge_stmt_1826_PhiAck/$entry
      -- CP-element group 344: 	 branch_block_stmt_1181/merge_stmt_1826_PhiAck/$exit
      -- CP-element group 344: 	 branch_block_stmt_1181/merge_stmt_1826_PhiAck/dummy
      -- 
    rr_4755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(344), ack => type_cast_1833_inst_req_0); -- 
    cr_4760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(344), ack => type_cast_1833_inst_req_1); -- 
    cr_4746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(344), ack => type_cast_1829_inst_req_1); -- 
    rr_4741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(344), ack => type_cast_1829_inst_req_0); -- 
    cr_4774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(344), ack => type_cast_1837_inst_req_1); -- 
    rr_4769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(344), ack => type_cast_1837_inst_req_0); -- 
    convolution3D_CP_3515_elements(344) <= OrReduce(convolution3D_CP_3515_elements(146) & convolution3D_CP_3515_elements(129));
    -- CP-element group 345:  transition  output  delay-element  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	166 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	349 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- CP-element group 345: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1951/$exit
      -- CP-element group 345: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/$exit
      -- CP-element group 345: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1955_konst_delay_trans
      -- CP-element group 345: 	 branch_block_stmt_1181/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_req
      -- 
    phi_stmt_1951_req_6246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1951_req_6246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(345), ack => phi_stmt_1951_req_0); -- 
    -- Element group convolution3D_CP_3515_elements(345) is a control-delay.
    cp_element_345_delay: control_delay_element  generic map(name => " 345_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(166), ack => convolution3D_CP_3515_elements(345), clk => clk, reset =>reset);
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	208 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (2) 
      -- CP-element group 346: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/Sample/ra
      -- 
    ra_6266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_0, ack => convolution3D_CP_3515_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	208 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (2) 
      -- CP-element group 347: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/Update/ca
      -- 
    ca_6271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_1, ack => convolution3D_CP_3515_elements(347)); -- 
    -- CP-element group 348:  join  transition  output  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	349 
    -- CP-element group 348:  members (6) 
      -- CP-element group 348: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- CP-element group 348: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/$exit
      -- CP-element group 348: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/$exit
      -- CP-element group 348: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/$exit
      -- CP-element group 348: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_sources/type_cast_1957/SplitProtocol/$exit
      -- CP-element group 348: 	 branch_block_stmt_1181/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1951/phi_stmt_1951_req
      -- 
    phi_stmt_1951_req_6272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1951_req_6272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(348), ack => phi_stmt_1951_req_1); -- 
    convolution3D_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(346) & convolution3D_CP_3515_elements(347);
      gj_convolution3D_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  merge  transition  place  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	345 
    -- CP-element group 349: 	348 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (2) 
      -- CP-element group 349: 	 branch_block_stmt_1181/merge_stmt_1950_PhiReqMerge
      -- CP-element group 349: 	 branch_block_stmt_1181/merge_stmt_1950_PhiAck/$entry
      -- 
    convolution3D_CP_3515_elements(349) <= OrReduce(convolution3D_CP_3515_elements(345) & convolution3D_CP_3515_elements(348));
    -- CP-element group 350:  fork  transition  place  input  output  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	198 
    -- CP-element group 350: 	186 
    -- CP-element group 350: 	205 
    -- CP-element group 350: 	202 
    -- CP-element group 350: 	194 
    -- CP-element group 350: 	174 
    -- CP-element group 350: 	182 
    -- CP-element group 350: 	190 
    -- CP-element group 350: 	167 
    -- CP-element group 350: 	168 
    -- CP-element group 350: 	170 
    -- CP-element group 350: 	171 
    -- CP-element group 350: 	178 
    -- CP-element group 350:  members (56) 
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_resized_1
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_Update/req
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_scale_1/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_resize_1/index_resize_ack
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_update_start
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113__entry__
      -- CP-element group 350: 	 branch_block_stmt_1181/merge_stmt_1950__exit__
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_scale_1/$exit
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_resize_1/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_resize_1/index_resize_req
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_sample_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_resize_1/$exit
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/addr_of_1964_complete/req
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_scale_1/scale_rename_req
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_scale_1/scale_rename_ack
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_computed_1
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_index_scaled_1
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/array_obj_ref_1963_final_index_sum_regn_Sample/req
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_Sample/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/RPIPE_maxpool_input_pipe_1967_Sample/rr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1971_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_1984_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2002_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2020_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2038_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2056_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2074_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/type_cast_2092_Update/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Update/word_access_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Update/word_access_complete/word_0/$entry
      -- CP-element group 350: 	 branch_block_stmt_1181/assign_stmt_1965_to_assign_stmt_2113/ptr_deref_2100_Update/word_access_complete/word_0/cr
      -- CP-element group 350: 	 branch_block_stmt_1181/merge_stmt_1950_PhiAck/$exit
      -- CP-element group 350: 	 branch_block_stmt_1181/merge_stmt_1950_PhiAck/phi_stmt_1951_ack
      -- 
    phi_stmt_1951_ack_6277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1951_ack_0, ack => convolution3D_CP_3515_elements(350)); -- 
    req_4900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => array_obj_ref_1963_index_offset_req_1); -- 
    req_4915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => addr_of_1964_final_reg_req_1); -- 
    req_4895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => array_obj_ref_1963_index_offset_req_0); -- 
    rr_4924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => RPIPE_maxpool_input_pipe_1967_inst_req_0); -- 
    cr_4943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => type_cast_1971_inst_req_1); -- 
    cr_4971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => type_cast_1984_inst_req_1); -- 
    cr_4999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => type_cast_2002_inst_req_1); -- 
    cr_5027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => type_cast_2020_inst_req_1); -- 
    cr_5055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => type_cast_2038_inst_req_1); -- 
    cr_5083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => type_cast_2056_inst_req_1); -- 
    cr_5111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => type_cast_2074_inst_req_1); -- 
    cr_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => type_cast_2092_inst_req_1); -- 
    cr_5189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(350), ack => ptr_deref_2100_store_0_req_1); -- 
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	207 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (2) 
      -- CP-element group 351: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/Sample/ra
      -- 
    ra_6309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2151_inst_ack_0, ack => convolution3D_CP_3515_elements(351)); -- 
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	207 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (2) 
      -- CP-element group 352: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/Update/ca
      -- 
    ca_6314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2151_inst_ack_1, ack => convolution3D_CP_3515_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (6) 
      -- CP-element group 353: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- CP-element group 353: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/$exit
      -- CP-element group 353: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/$exit
      -- CP-element group 353: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/$exit
      -- CP-element group 353: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2151/SplitProtocol/$exit
      -- CP-element group 353: 	 branch_block_stmt_1181/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_req
      -- 
    phi_stmt_2145_req_6315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2145_req_6315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(353), ack => phi_stmt_2145_req_1); -- 
    convolution3D_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(351) & convolution3D_CP_3515_elements(352);
      gj_convolution3D_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  transition  output  delay-element  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	155 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (5) 
      -- CP-element group 354: 	 branch_block_stmt_1181/ifx_xend_forx_xend215_PhiReq/$exit
      -- CP-element group 354: 	 branch_block_stmt_1181/ifx_xend_forx_xend215_PhiReq/phi_stmt_2145/$exit
      -- CP-element group 354: 	 branch_block_stmt_1181/ifx_xend_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/$exit
      -- CP-element group 354: 	 branch_block_stmt_1181/ifx_xend_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_sources/type_cast_2149_konst_delay_trans
      -- CP-element group 354: 	 branch_block_stmt_1181/ifx_xend_forx_xend215_PhiReq/phi_stmt_2145/phi_stmt_2145_req
      -- 
    phi_stmt_2145_req_6326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2145_req_6326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(354), ack => phi_stmt_2145_req_0); -- 
    -- Element group convolution3D_CP_3515_elements(354) is a control-delay.
    cp_element_354_delay: control_delay_element  generic map(name => " 354_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(155), ack => convolution3D_CP_3515_elements(354), clk => clk, reset =>reset);
    -- CP-element group 355:  merge  transition  place  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (2) 
      -- CP-element group 355: 	 branch_block_stmt_1181/merge_stmt_2144_PhiReqMerge
      -- CP-element group 355: 	 branch_block_stmt_1181/merge_stmt_2144_PhiAck/$entry
      -- 
    convolution3D_CP_3515_elements(355) <= OrReduce(convolution3D_CP_3515_elements(353) & convolution3D_CP_3515_elements(354));
    -- CP-element group 356:  branch  transition  place  input  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	209 
    -- CP-element group 356: 	210 
    -- CP-element group 356:  members (15) 
      -- CP-element group 356: 	 branch_block_stmt_1181/assign_stmt_2158_to_assign_stmt_2164__entry__
      -- CP-element group 356: 	 branch_block_stmt_1181/merge_stmt_2144__exit__
      -- CP-element group 356: 	 branch_block_stmt_1181/if_stmt_2165__entry__
      -- CP-element group 356: 	 branch_block_stmt_1181/assign_stmt_2158_to_assign_stmt_2164__exit__
      -- CP-element group 356: 	 branch_block_stmt_1181/assign_stmt_2158_to_assign_stmt_2164/$entry
      -- CP-element group 356: 	 branch_block_stmt_1181/assign_stmt_2158_to_assign_stmt_2164/$exit
      -- CP-element group 356: 	 branch_block_stmt_1181/if_stmt_2165_dead_link/$entry
      -- CP-element group 356: 	 branch_block_stmt_1181/if_stmt_2165_eval_test/$entry
      -- CP-element group 356: 	 branch_block_stmt_1181/if_stmt_2165_eval_test/$exit
      -- CP-element group 356: 	 branch_block_stmt_1181/if_stmt_2165_eval_test/branch_req
      -- CP-element group 356: 	 branch_block_stmt_1181/R_tobool218_2166_place
      -- CP-element group 356: 	 branch_block_stmt_1181/if_stmt_2165_if_link/$entry
      -- CP-element group 356: 	 branch_block_stmt_1181/if_stmt_2165_else_link/$entry
      -- CP-element group 356: 	 branch_block_stmt_1181/merge_stmt_2144_PhiAck/$exit
      -- CP-element group 356: 	 branch_block_stmt_1181/merge_stmt_2144_PhiAck/phi_stmt_2145_ack
      -- 
    phi_stmt_2145_ack_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2145_ack_0, ack => convolution3D_CP_3515_elements(356)); -- 
    branch_req_5223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(356), ack => if_stmt_2165_branch_req_0); -- 
    -- CP-element group 357:  transition  output  delay-element  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	212 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (4) 
      -- CP-element group 357: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/$exit
      -- CP-element group 357: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/$exit
      -- CP-element group 357: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2203_konst_delay_trans
      -- CP-element group 357: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_req
      -- 
    phi_stmt_2197_req_6354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2197_req_6354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(357), ack => phi_stmt_2197_req_1); -- 
    -- Element group convolution3D_CP_3515_elements(357) is a control-delay.
    cp_element_357_delay: control_delay_element  generic map(name => " 357_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(212), ack => convolution3D_CP_3515_elements(357), clk => clk, reset =>reset);
    -- CP-element group 358:  transition  output  delay-element  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	212 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (4) 
      -- CP-element group 358: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/$exit
      -- CP-element group 358: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$exit
      -- CP-element group 358: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2196_konst_delay_trans
      -- CP-element group 358: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_req
      -- 
    phi_stmt_2190_req_6362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2190_req_6362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(358), ack => phi_stmt_2190_req_1); -- 
    -- Element group convolution3D_CP_3515_elements(358) is a control-delay.
    cp_element_358_delay: control_delay_element  generic map(name => " 358_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(212), ack => convolution3D_CP_3515_elements(358), clk => clk, reset =>reset);
    -- CP-element group 359:  join  transition  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	367 
    -- CP-element group 359:  members (1) 
      -- CP-element group 359: 	 branch_block_stmt_1181/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(358) & convolution3D_CP_3515_elements(357);
      gj_convolution3D_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	220 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	362 
    -- CP-element group 360:  members (2) 
      -- CP-element group 360: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/Sample/ra
      -- 
    ra_6382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2200_inst_ack_0, ack => convolution3D_CP_3515_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	220 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (2) 
      -- CP-element group 361: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/Update/ca
      -- 
    ca_6387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2200_inst_ack_1, ack => convolution3D_CP_3515_elements(361)); -- 
    -- CP-element group 362:  join  transition  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	366 
    -- CP-element group 362:  members (5) 
      -- CP-element group 362: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/$exit
      -- CP-element group 362: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/$exit
      -- CP-element group 362: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/$exit
      -- CP-element group 362: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_sources/type_cast_2200/SplitProtocol/$exit
      -- CP-element group 362: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2197/phi_stmt_2197_req
      -- 
    phi_stmt_2197_req_6388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2197_req_6388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(362), ack => phi_stmt_2197_req_0); -- 
    convolution3D_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(360) & convolution3D_CP_3515_elements(361);
      gj_convolution3D_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	220 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	365 
    -- CP-element group 363:  members (2) 
      -- CP-element group 363: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Sample/ra
      -- 
    ra_6405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_0, ack => convolution3D_CP_3515_elements(363)); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	220 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (2) 
      -- CP-element group 364: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/Update/ca
      -- 
    ca_6410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2193_inst_ack_1, ack => convolution3D_CP_3515_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (5) 
      -- CP-element group 365: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/$exit
      -- CP-element group 365: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/$exit
      -- CP-element group 365: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/$exit
      -- CP-element group 365: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_sources/type_cast_2193/SplitProtocol/$exit
      -- CP-element group 365: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_2190/phi_stmt_2190_req
      -- 
    phi_stmt_2190_req_6411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2190_req_6411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(365), ack => phi_stmt_2190_req_0); -- 
    convolution3D_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(363) & convolution3D_CP_3515_elements(364);
      gj_convolution3D_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	362 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (1) 
      -- CP-element group 366: 	 branch_block_stmt_1181/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(362) & convolution3D_CP_3515_elements(365);
      gj_convolution3D_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  merge  fork  transition  place  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	359 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_1181/merge_stmt_2189_PhiReqMerge
      -- CP-element group 367: 	 branch_block_stmt_1181/merge_stmt_2189_PhiAck/$entry
      -- 
    convolution3D_CP_3515_elements(367) <= OrReduce(convolution3D_CP_3515_elements(359) & convolution3D_CP_3515_elements(366));
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (1) 
      -- CP-element group 368: 	 branch_block_stmt_1181/merge_stmt_2189_PhiAck/phi_stmt_2190_ack
      -- 
    phi_stmt_2190_ack_6416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2190_ack_0, ack => convolution3D_CP_3515_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (1) 
      -- CP-element group 369: 	 branch_block_stmt_1181/merge_stmt_2189_PhiAck/phi_stmt_2197_ack
      -- 
    phi_stmt_2197_ack_6417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2197_ack_0, ack => convolution3D_CP_3515_elements(369)); -- 
    -- CP-element group 370:  join  fork  transition  place  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	217 
    -- CP-element group 370: 	218 
    -- CP-element group 370: 	213 
    -- CP-element group 370: 	216 
    -- CP-element group 370:  members (16) 
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243__entry__
      -- CP-element group 370: 	 branch_block_stmt_1181/merge_stmt_2189__exit__
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/$entry
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/RPIPE_maxpool_input_pipe_2218_Sample/rr
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_update_start_
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2222_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_update_start_
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_Sample/rr
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_1181/assign_stmt_2210_to_assign_stmt_2243/type_cast_2237_Update/cr
      -- CP-element group 370: 	 branch_block_stmt_1181/merge_stmt_2189_PhiAck/$exit
      -- 
    rr_5262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(370), ack => RPIPE_maxpool_input_pipe_2218_inst_req_0); -- 
    cr_5281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(370), ack => type_cast_2222_inst_req_1); -- 
    rr_5290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(370), ack => type_cast_2237_inst_req_0); -- 
    cr_5295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(370), ack => type_cast_2237_inst_req_1); -- 
    convolution3D_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(368) & convolution3D_CP_3515_elements(369);
      gj_convolution3D_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	221 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	373 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Sample/ra
      -- 
    ra_6441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2254_inst_ack_0, ack => convolution3D_CP_3515_elements(371)); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	221 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (2) 
      -- CP-element group 372: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/Update/ca
      -- 
    ca_6446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2254_inst_ack_1, ack => convolution3D_CP_3515_elements(372)); -- 
    -- CP-element group 373:  join  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	371 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (8) 
      -- CP-element group 373: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/$exit
      -- CP-element group 373: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/$exit
      -- CP-element group 373: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/$exit
      -- CP-element group 373: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/$exit
      -- CP-element group 373: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_sources/type_cast_2254/SplitProtocol/$exit
      -- CP-element group 373: 	 branch_block_stmt_1181/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_2251/phi_stmt_2251_req
      -- CP-element group 373: 	 branch_block_stmt_1181/merge_stmt_2250_PhiReqMerge
      -- CP-element group 373: 	 branch_block_stmt_1181/merge_stmt_2250_PhiAck/$entry
      -- 
    phi_stmt_2251_req_6447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2251_req_6447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(373), ack => phi_stmt_2251_req_0); -- 
    convolution3D_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(371) & convolution3D_CP_3515_elements(372);
      gj_convolution3D_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	222 
    -- CP-element group 374: 	223 
    -- CP-element group 374: 	225 
    -- CP-element group 374: 	227 
    -- CP-element group 374:  members (29) 
      -- CP-element group 374: 	 branch_block_stmt_1181/merge_stmt_2250__exit__
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289__entry__
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_update_start_
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_resized_1
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_scaled_1
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_computed_1
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_resize_1/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_resize_1/$exit
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_resize_1/index_resize_req
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_resize_1/index_resize_ack
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_scale_1/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_scale_1/$exit
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_scale_1/scale_rename_req
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_index_scale_1/scale_rename_ack
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_update_start
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_Sample/req
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/array_obj_ref_2283_final_index_sum_regn_Update/req
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_complete/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/addr_of_2284_complete/req
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_update_start_
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Update/word_access_complete/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Update/word_access_complete/word_0/$entry
      -- CP-element group 374: 	 branch_block_stmt_1181/assign_stmt_2261_to_assign_stmt_2289/ptr_deref_2287_Update/word_access_complete/word_0/cr
      -- CP-element group 374: 	 branch_block_stmt_1181/merge_stmt_2250_PhiAck/$exit
      -- CP-element group 374: 	 branch_block_stmt_1181/merge_stmt_2250_PhiAck/phi_stmt_2251_ack
      -- 
    phi_stmt_2251_ack_6452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2251_ack_0, ack => convolution3D_CP_3515_elements(374)); -- 
    req_5343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(374), ack => array_obj_ref_2283_index_offset_req_0); -- 
    req_5348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(374), ack => array_obj_ref_2283_index_offset_req_1); -- 
    req_5363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(374), ack => addr_of_2284_final_reg_req_1); -- 
    cr_5413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(374), ack => ptr_deref_2287_store_0_req_1); -- 
    -- CP-element group 375:  merge  place  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	228 
    -- CP-element group 375: 	209 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (1) 
      -- CP-element group 375: 	 branch_block_stmt_1181/merge_stmt_2291_PhiReqMerge
      -- 
    convolution3D_CP_3515_elements(375) <= OrReduce(convolution3D_CP_3515_elements(228) & convolution3D_CP_3515_elements(209));
    -- CP-element group 376:  join  fork  transition  place  output  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	229 
    -- CP-element group 376: 	230 
    -- CP-element group 376:  members (36) 
      -- CP-element group 376: 	 branch_block_stmt_1181/merge_stmt_2291__exit__
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304__entry__
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_word_addrgen/root_register_req
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_word_addrgen/root_register_ack
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Update/word_access_complete/word_0/cr
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Update/word_access_complete/word_0/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Update/word_access_complete/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_word_addrgen/$exit
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/word_access_start/word_0/rr
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/word_access_start/word_0/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/word_access_start/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/ptr_deref_2301_Split/split_ack
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/ptr_deref_2301_Split/split_req
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/ptr_deref_2301_Split/$exit
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_Sample/ptr_deref_2301_Split/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_word_addrgen/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_sample_start_
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_update_start_
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_word_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_root_address_calculated
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_address_resized
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_addr_resize/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_addr_resize/$exit
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_addr_resize/base_resize_req
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_addr_resize/base_resize_ack
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_plus_offset/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_plus_offset/$exit
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_plus_offset/sum_rename_req
      -- CP-element group 376: 	 branch_block_stmt_1181/assign_stmt_2299_to_assign_stmt_2304/ptr_deref_2301_base_plus_offset/sum_rename_ack
      -- CP-element group 376: 	 branch_block_stmt_1181/merge_stmt_2291_PhiAck/$entry
      -- CP-element group 376: 	 branch_block_stmt_1181/merge_stmt_2291_PhiAck/$exit
      -- CP-element group 376: 	 branch_block_stmt_1181/merge_stmt_2291_PhiAck/dummy
      -- 
    cr_5466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(376), ack => ptr_deref_2301_store_0_req_1); -- 
    rr_5455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(376), ack => ptr_deref_2301_store_0_req_0); -- 
    convolution3D_CP_3515_elements(376) <= convolution3D_CP_3515_elements(375);
    -- CP-element group 377:  transition  output  delay-element  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	244 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	381 
    -- CP-element group 377:  members (5) 
      -- CP-element group 377: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- CP-element group 377: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2350/$exit
      -- CP-element group 377: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/$exit
      -- CP-element group 377: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2354_konst_delay_trans
      -- CP-element group 377: 	 branch_block_stmt_1181/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_req
      -- 
    phi_stmt_2350_req_6474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2350_req_6474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(377), ack => phi_stmt_2350_req_0); -- 
    -- Element group convolution3D_CP_3515_elements(377) is a control-delay.
    cp_element_377_delay: control_delay_element  generic map(name => " 377_delay", delay_value => 1)  port map(req => convolution3D_CP_3515_elements(244), ack => convolution3D_CP_3515_elements(377), clk => clk, reset =>reset);
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	255 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378:  members (2) 
      -- CP-element group 378: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/Sample/ra
      -- 
    ra_6494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2356_inst_ack_0, ack => convolution3D_CP_3515_elements(378)); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	255 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (2) 
      -- CP-element group 379: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/Update/ca
      -- 
    ca_6499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2356_inst_ack_1, ack => convolution3D_CP_3515_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	381 
    -- CP-element group 380:  members (6) 
      -- CP-element group 380: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 380: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/$exit
      -- CP-element group 380: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/$exit
      -- CP-element group 380: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/$exit
      -- CP-element group 380: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_sources/type_cast_2356/SplitProtocol/$exit
      -- CP-element group 380: 	 branch_block_stmt_1181/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_2350/phi_stmt_2350_req
      -- 
    phi_stmt_2350_req_6500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2350_req_6500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(380), ack => phi_stmt_2350_req_1); -- 
    convolution3D_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_3515_elements(378) & convolution3D_CP_3515_elements(379);
      gj_convolution3D_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_3515_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  merge  transition  place  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	377 
    -- CP-element group 381: 	380 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (2) 
      -- CP-element group 381: 	 branch_block_stmt_1181/merge_stmt_2349_PhiReqMerge
      -- CP-element group 381: 	 branch_block_stmt_1181/merge_stmt_2349_PhiAck/$entry
      -- 
    convolution3D_CP_3515_elements(381) <= OrReduce(convolution3D_CP_3515_elements(377) & convolution3D_CP_3515_elements(380));
    -- CP-element group 382:  fork  transition  place  input  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	245 
    -- CP-element group 382: 	249 
    -- CP-element group 382: 	250 
    -- CP-element group 382: 	251 
    -- CP-element group 382: 	252 
    -- CP-element group 382:  members (20) 
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392__entry__
      -- CP-element group 382: 	 branch_block_stmt_1181/merge_stmt_2349__exit__
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_Sample/$entry
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_Sample/req
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_Sample/$entry
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/WPIPE_num_out_pipe_2363_sample_start_
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/$entry
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_update_start_
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_sample_start_
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_Update/ccr
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_Sample/crr
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_Sample/$entry
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_update_start_
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2377_sample_start_
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_Update/ccr
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_1181/assign_stmt_2362_to_assign_stmt_2392/call_stmt_2381_Sample/crr
      -- CP-element group 382: 	 branch_block_stmt_1181/merge_stmt_2349_PhiAck/$exit
      -- CP-element group 382: 	 branch_block_stmt_1181/merge_stmt_2349_PhiAck/phi_stmt_2350_ack
      -- 
    phi_stmt_2350_ack_6505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2350_ack_0, ack => convolution3D_CP_3515_elements(382)); -- 
    req_5568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(382), ack => WPIPE_num_out_pipe_2363_inst_req_0); -- 
    ccr_5601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(382), ack => call_stmt_2377_call_req_1); -- 
    crr_5596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(382), ack => call_stmt_2377_call_req_0); -- 
    ccr_5615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_5615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(382), ack => call_stmt_2381_call_req_1); -- 
    crr_5610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_5610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_3515_elements(382), ack => call_stmt_2381_call_req_0); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1679_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1866_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_2140_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_2455_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1796 : std_logic_vector(63 downto 0);
    signal R_indvar411_1962_resized : std_logic_vector(13 downto 0);
    signal R_indvar411_1962_scaled : std_logic_vector(13 downto 0);
    signal R_indvar425_1501_resized : std_logic_vector(13 downto 0);
    signal R_indvar425_1501_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1817_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1817_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_2282_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_2282_scaled : std_logic_vector(13 downto 0);
    signal add102_1547 : std_logic_vector(63 downto 0);
    signal add108_1565 : std_logic_vector(63 downto 0);
    signal add114_1583 : std_logic_vector(63 downto 0);
    signal add120_1601 : std_logic_vector(63 downto 0);
    signal add1216x_xi370_2267 : std_logic_vector(63 downto 0);
    signal add1216x_xi_1802 : std_logic_vector(63 downto 0);
    signal add126_1619 : std_logic_vector(63 downto 0);
    signal add132_1637 : std_logic_vector(63 downto 0);
    signal add13_1232 : std_logic_vector(15 downto 0);
    signal add171_1990 : std_logic_vector(63 downto 0);
    signal add177_2008 : std_logic_vector(63 downto 0);
    signal add183_2026 : std_logic_vector(63 downto 0);
    signal add189_2044 : std_logic_vector(63 downto 0);
    signal add195_2062 : std_logic_vector(63 downto 0);
    signal add201_2080 : std_logic_vector(63 downto 0);
    signal add207_2098 : std_logic_vector(63 downto 0);
    signal add23_1257 : std_logic_vector(15 downto 0);
    signal add33_1282 : std_logic_vector(15 downto 0);
    signal add43_1307 : std_logic_vector(15 downto 0);
    signal add53_1332 : std_logic_vector(15 downto 0);
    signal add63_1357 : std_logic_vector(63 downto 0);
    signal add73_1382 : std_logic_vector(15 downto 0);
    signal add96_1529 : std_logic_vector(63 downto 0);
    signal add_1207 : std_logic_vector(31 downto 0);
    signal addx_xi361_2228 : std_logic_vector(63 downto 0);
    signal addx_xi_1763 : std_logic_vector(63 downto 0);
    signal and217_2158 : std_logic_vector(63 downto 0);
    signal and_1697 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1502_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1502_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1502_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1502_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1502_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1502_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1818_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1818_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1818_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1818_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1818_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1818_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1963_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1963_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1963_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1963_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1963_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1963_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2283_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2283_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2283_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2283_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2283_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2283_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_1820 : std_logic_vector(31 downto 0);
    signal arrayidx211_1965 : std_logic_vector(31 downto 0);
    signal arrayidx226_2285 : std_logic_vector(31 downto 0);
    signal arrayidx_1504 : std_logic_vector(31 downto 0);
    signal call105_1556 : std_logic_vector(7 downto 0);
    signal call111_1574 : std_logic_vector(7 downto 0);
    signal call117_1592 : std_logic_vector(7 downto 0);
    signal call11_1223 : std_logic_vector(7 downto 0);
    signal call123_1610 : std_logic_vector(7 downto 0);
    signal call129_1628 : std_logic_vector(7 downto 0);
    signal call164_1968 : std_logic_vector(7 downto 0);
    signal call168_1981 : std_logic_vector(7 downto 0);
    signal call16_1235 : std_logic_vector(7 downto 0);
    signal call174_1999 : std_logic_vector(7 downto 0);
    signal call180_2017 : std_logic_vector(7 downto 0);
    signal call186_2035 : std_logic_vector(7 downto 0);
    signal call192_2053 : std_logic_vector(7 downto 0);
    signal call198_2071 : std_logic_vector(7 downto 0);
    signal call204_2089 : std_logic_vector(7 downto 0);
    signal call21_1248 : std_logic_vector(7 downto 0);
    signal call229_2307 : std_logic_vector(63 downto 0);
    signal call26_1260 : std_logic_vector(7 downto 0);
    signal call270_2407 : std_logic_vector(7 downto 0);
    signal call273_2411 : std_logic_vector(7 downto 0);
    signal call275_2414 : std_logic_vector(63 downto 0);
    signal call2_1198 : std_logic_vector(7 downto 0);
    signal call31_1273 : std_logic_vector(7 downto 0);
    signal call36_1285 : std_logic_vector(7 downto 0);
    signal call41_1298 : std_logic_vector(7 downto 0);
    signal call46_1310 : std_logic_vector(7 downto 0);
    signal call51_1323 : std_logic_vector(7 downto 0);
    signal call56_1335 : std_logic_vector(7 downto 0);
    signal call61_1348 : std_logic_vector(7 downto 0);
    signal call66_1360 : std_logic_vector(7 downto 0);
    signal call6_1210 : std_logic_vector(7 downto 0);
    signal call71_1373 : std_logic_vector(7 downto 0);
    signal call89_1507 : std_logic_vector(7 downto 0);
    signal call93_1520 : std_logic_vector(7 downto 0);
    signal call99_1538 : std_logic_vector(7 downto 0);
    signal call_1185 : std_logic_vector(7 downto 0);
    signal callx_xi359_2219 : std_logic_vector(7 downto 0);
    signal callx_xi_1754 : std_logic_vector(7 downto 0);
    signal cmp161379_1874 : std_logic_vector(0 downto 0);
    signal cmp383_1411 : std_logic_vector(0 downto 0);
    signal cmpx_xi364_2243 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1778 : std_logic_vector(0 downto 0);
    signal conv101_1542 : std_logic_vector(63 downto 0);
    signal conv107_1560 : std_logic_vector(63 downto 0);
    signal conv113_1578 : std_logic_vector(63 downto 0);
    signal conv119_1596 : std_logic_vector(63 downto 0);
    signal conv125_1614 : std_logic_vector(63 downto 0);
    signal conv12_1227 : std_logic_vector(15 downto 0);
    signal conv131_1632 : std_logic_vector(63 downto 0);
    signal conv145_1830 : std_logic_vector(63 downto 0);
    signal conv147_1834 : std_logic_vector(63 downto 0);
    signal conv153_1838 : std_logic_vector(63 downto 0);
    signal conv155_1868 : std_logic_vector(63 downto 0);
    signal conv165_1972 : std_logic_vector(63 downto 0);
    signal conv170_1985 : std_logic_vector(63 downto 0);
    signal conv176_2003 : std_logic_vector(63 downto 0);
    signal conv182_2021 : std_logic_vector(63 downto 0);
    signal conv188_2039 : std_logic_vector(63 downto 0);
    signal conv194_2057 : std_logic_vector(63 downto 0);
    signal conv19_1239 : std_logic_vector(15 downto 0);
    signal conv1_1189 : std_logic_vector(31 downto 0);
    signal conv200_2075 : std_logic_vector(63 downto 0);
    signal conv206_2093 : std_logic_vector(63 downto 0);
    signal conv22_1252 : std_logic_vector(15 downto 0);
    signal conv230_2404 : std_logic_vector(63 downto 0);
    signal conv254_2374 : std_logic_vector(63 downto 0);
    signal conv276_2419 : std_logic_vector(63 downto 0);
    signal conv281_2428 : std_logic_vector(63 downto 0);
    signal conv283_2432 : std_logic_vector(63 downto 0);
    signal conv288_2457 : std_logic_vector(63 downto 0);
    signal conv292_2464 : std_logic_vector(7 downto 0);
    signal conv298_2474 : std_logic_vector(7 downto 0);
    signal conv29_1264 : std_logic_vector(15 downto 0);
    signal conv2x_xi354_2181 : std_logic_vector(31 downto 0);
    signal conv2x_xi_1716 : std_logic_vector(31 downto 0);
    signal conv304_2484 : std_logic_vector(7 downto 0);
    signal conv310_2494 : std_logic_vector(7 downto 0);
    signal conv316_2504 : std_logic_vector(7 downto 0);
    signal conv322_2514 : std_logic_vector(7 downto 0);
    signal conv328_2524 : std_logic_vector(7 downto 0);
    signal conv32_1277 : std_logic_vector(15 downto 0);
    signal conv334_2534 : std_logic_vector(7 downto 0);
    signal conv39_1289 : std_logic_vector(15 downto 0);
    signal conv3_1202 : std_logic_vector(31 downto 0);
    signal conv42_1302 : std_logic_vector(15 downto 0);
    signal conv49_1314 : std_logic_vector(15 downto 0);
    signal conv52_1327 : std_logic_vector(15 downto 0);
    signal conv59_1339 : std_logic_vector(63 downto 0);
    signal conv5x_xi360_2223 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1758 : std_logic_vector(63 downto 0);
    signal conv62_1352 : std_logic_vector(63 downto 0);
    signal conv69_1364 : std_logic_vector(15 downto 0);
    signal conv72_1377 : std_logic_vector(15 downto 0);
    signal conv79_1386 : std_logic_vector(31 downto 0);
    signal conv81_1390 : std_logic_vector(31 downto 0);
    signal conv83_1405 : std_logic_vector(63 downto 0);
    signal conv90_1511 : std_logic_vector(63 downto 0);
    signal conv95_1524 : std_logic_vector(63 downto 0);
    signal conv9_1214 : std_logic_vector(15 downto 0);
    signal convx_xi363_2238 : std_logic_vector(31 downto 0);
    signal convx_xi_1773 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi358_2197 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_1732 : std_logic_vector(63 downto 0);
    signal exitcond28_1652 : std_logic_vector(0 downto 0);
    signal exitcond5_2392 : std_logic_vector(0 downto 0);
    signal exitcond_2113 : std_logic_vector(0 downto 0);
    signal iNsTr_35_1751 : std_logic_vector(15 downto 0);
    signal iNsTr_48_2299 : std_logic_vector(31 downto 0);
    signal iNsTr_59_2177 : std_logic_vector(63 downto 0);
    signal iNsTr_71_2216 : std_logic_vector(15 downto 0);
    signal iNsTr_97_2261 : std_logic_vector(63 downto 0);
    signal indvar411_1951 : std_logic_vector(63 downto 0);
    signal indvar425_1490 : std_logic_vector(63 downto 0);
    signal indvar_2350 : std_logic_vector(63 downto 0);
    signal indvarx_xnext412_2108 : std_logic_vector(63 downto 0);
    signal indvarx_xnext426_1647 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_2387 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_1684 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_2145 : std_logic_vector(63 downto 0);
    signal mul148_1843 : std_logic_vector(63 downto 0);
    signal mul151_1848 : std_logic_vector(63 downto 0);
    signal mul154_1853 : std_logic_vector(63 downto 0);
    signal mul253_2362 : std_logic_vector(63 downto 0);
    signal mul284_2438 : std_logic_vector(63 downto 0);
    signal mul287_2443 : std_logic_vector(63 downto 0);
    signal mul82_1400 : std_logic_vector(31 downto 0);
    signal mul_1395 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi357_2190 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_1725 : std_logic_vector(15 downto 0);
    signal phitmp387_2142 : std_logic_vector(63 downto 0);
    signal phitmp_1681 : std_logic_vector(63 downto 0);
    signal ptr_deref_1639_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1639_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1639_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1639_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1639_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1639_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1822_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1822_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1822_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1822_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1822_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1822_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2100_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2100_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2287_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2287_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2287_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2287_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2287_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2287_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2301_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2301_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2301_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2301_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2301_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2301_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext352_2448 : std_logic_vector(63 downto 0);
    signal sext_1859 : std_logic_vector(63 downto 0);
    signal sh_promx_xi371_2273 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1808 : std_logic_vector(63 downto 0);
    signal shl104_1553 : std_logic_vector(63 downto 0);
    signal shl10_1220 : std_logic_vector(15 downto 0);
    signal shl110_1571 : std_logic_vector(63 downto 0);
    signal shl116_1589 : std_logic_vector(63 downto 0);
    signal shl122_1607 : std_logic_vector(63 downto 0);
    signal shl128_1625 : std_logic_vector(63 downto 0);
    signal shl14x_xi372_2278 : std_logic_vector(63 downto 0);
    signal shl14x_xi_1813 : std_logic_vector(63 downto 0);
    signal shl167_1978 : std_logic_vector(63 downto 0);
    signal shl173_1996 : std_logic_vector(63 downto 0);
    signal shl179_2014 : std_logic_vector(63 downto 0);
    signal shl185_2032 : std_logic_vector(63 downto 0);
    signal shl191_2050 : std_logic_vector(63 downto 0);
    signal shl197_2068 : std_logic_vector(63 downto 0);
    signal shl203_2086 : std_logic_vector(63 downto 0);
    signal shl20_1245 : std_logic_vector(15 downto 0);
    signal shl30_1270 : std_logic_vector(15 downto 0);
    signal shl40_1295 : std_logic_vector(15 downto 0);
    signal shl50_1320 : std_logic_vector(15 downto 0);
    signal shl60_1345 : std_logic_vector(63 downto 0);
    signal shl70_1370 : std_logic_vector(15 downto 0);
    signal shl8x_xi362_2234 : std_logic_vector(63 downto 0);
    signal shl8x_xi362x_xlcssa_2251 : std_logic_vector(63 downto 0);
    signal shl8x_xi_1769 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_1786 : std_logic_vector(63 downto 0);
    signal shl92_1517 : std_logic_vector(63 downto 0);
    signal shl98_1535 : std_logic_vector(63 downto 0);
    signal shl_1195 : std_logic_vector(31 downto 0);
    signal shlx_xi355_2187 : std_logic_vector(31 downto 0);
    signal shlx_xi_1722 : std_logic_vector(31 downto 0);
    signal shr295_2470 : std_logic_vector(63 downto 0);
    signal shr301_2480 : std_logic_vector(63 downto 0);
    signal shr307_2490 : std_logic_vector(63 downto 0);
    signal shr313_2500 : std_logic_vector(63 downto 0);
    signal shr319_2510 : std_logic_vector(63 downto 0);
    signal shr325_2520 : std_logic_vector(63 downto 0);
    signal shr331_2530 : std_logic_vector(63 downto 0);
    signal sub_2424 : std_logic_vector(63 downto 0);
    signal tmp10_1902 : std_logic_vector(63 downto 0);
    signal tmp11_1906 : std_logic_vector(63 downto 0);
    signal tmp12_1911 : std_logic_vector(63 downto 0);
    signal tmp13_1915 : std_logic_vector(63 downto 0);
    signal tmp14_1920 : std_logic_vector(63 downto 0);
    signal tmp15_1924 : std_logic_vector(31 downto 0);
    signal tmp16_1929 : std_logic_vector(63 downto 0);
    signal tmp17_1935 : std_logic_vector(63 downto 0);
    signal tmp18_1941 : std_logic_vector(0 downto 0);
    signal tmp20_1449 : std_logic_vector(31 downto 0);
    signal tmp21_1454 : std_logic_vector(31 downto 0);
    signal tmp22_1458 : std_logic_vector(31 downto 0);
    signal tmp23_1463 : std_logic_vector(31 downto 0);
    signal tmp24_1468 : std_logic_vector(63 downto 0);
    signal tmp25_1474 : std_logic_vector(63 downto 0);
    signal tmp26_1480 : std_logic_vector(0 downto 0);
    signal tmp388_2210 : std_logic_vector(15 downto 0);
    signal tmp389_2323 : std_logic_vector(15 downto 0);
    signal tmp393_2328 : std_logic_vector(15 downto 0);
    signal tmp3_2332 : std_logic_vector(63 downto 0);
    signal tmp406_1887 : std_logic_vector(63 downto 0);
    signal tmp407_1893 : std_logic_vector(0 downto 0);
    signal tmp408_2133 : std_logic_vector(63 downto 0);
    signal tmp415_1423 : std_logic_vector(31 downto 0);
    signal tmp417_1428 : std_logic_vector(31 downto 0);
    signal tmp418_1433 : std_logic_vector(63 downto 0);
    signal tmp419_1439 : std_logic_vector(63 downto 0);
    signal tmp420_1445 : std_logic_vector(0 downto 0);
    signal tmp422_1672 : std_logic_vector(63 downto 0);
    signal tmp4_2338 : std_logic_vector(63 downto 0);
    signal tmp6_2342 : std_logic_vector(63 downto 0);
    signal tmp7_2347 : std_logic_vector(63 downto 0);
    signal tmp9_1897 : std_logic_vector(63 downto 0);
    signal tmp_1745 : std_logic_vector(15 downto 0);
    signal tobool218_2164 : std_logic_vector(0 downto 0);
    signal tobool_1703 : std_logic_vector(0 downto 0);
    signal type_cast_1193_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1218_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1243_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1293_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1318_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1343_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1368_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1403_wire : std_logic_vector(63 downto 0);
    signal type_cast_1409_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1431_wire : std_logic_vector(63 downto 0);
    signal type_cast_1437_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1443_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1466_wire : std_logic_vector(63 downto 0);
    signal type_cast_1472_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1478_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1485_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1493_wire : std_logic_vector(63 downto 0);
    signal type_cast_1496_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1515_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1533_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1551_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1569_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1587_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1605_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1623_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1645_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1664_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1670_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1675_wire : std_logic_vector(63 downto 0);
    signal type_cast_1678_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1687_wire : std_logic_vector(63 downto 0);
    signal type_cast_1690_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1695_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1714_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1720_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1729_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1731_wire : std_logic_vector(15 downto 0);
    signal type_cast_1736_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1738_wire : std_logic_vector(63 downto 0);
    signal type_cast_1743_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1749_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1767_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1789_wire : std_logic_vector(63 downto 0);
    signal type_cast_1794_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1800_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1806_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1857_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1862_wire : std_logic_vector(63 downto 0);
    signal type_cast_1865_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1872_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1885_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1891_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1927_wire : std_logic_vector(63 downto 0);
    signal type_cast_1933_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1939_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1946_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1955_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1957_wire : std_logic_vector(63 downto 0);
    signal type_cast_1976_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1994_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2012_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2030_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2048_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2066_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2084_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2106_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2125_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2131_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2136_wire : std_logic_vector(63 downto 0);
    signal type_cast_2139_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2149_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2151_wire : std_logic_vector(63 downto 0);
    signal type_cast_2156_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2162_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2175_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2185_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2193_wire : std_logic_vector(15 downto 0);
    signal type_cast_2196_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2200_wire : std_logic_vector(63 downto 0);
    signal type_cast_2203_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2208_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2214_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2232_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2254_wire : std_logic_vector(63 downto 0);
    signal type_cast_2259_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2265_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2271_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2303_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2321_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2336_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2354_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2356_wire : std_logic_vector(63 downto 0);
    signal type_cast_2372_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2385_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2402_wire : std_logic_vector(63 downto 0);
    signal type_cast_2417_wire : std_logic_vector(63 downto 0);
    signal type_cast_2436_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2451_wire : std_logic_vector(63 downto 0);
    signal type_cast_2454_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2468_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2478_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2488_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2498_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2508_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2518_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2528_wire_constant : std_logic_vector(63 downto 0);
    signal umax19_1948 : std_logic_vector(63 downto 0);
    signal umax27_1487 : std_logic_vector(63 downto 0);
    signal umax421_1666 : std_logic_vector(63 downto 0);
    signal umax_2127 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1502_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1502_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1502_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1502_resized_base_address <= "00000000000000";
    array_obj_ref_1818_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1818_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1818_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1818_resized_base_address <= "00000000000000";
    array_obj_ref_1963_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1963_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1963_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1963_resized_base_address <= "00000000000000";
    array_obj_ref_2283_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2283_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2283_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2283_resized_base_address <= "00000000000000";
    iNsTr_48_2299 <= "00000000000000000000000000000000";
    ptr_deref_1639_word_offset_0 <= "00000000000000";
    ptr_deref_1822_word_offset_0 <= "00000000000000";
    ptr_deref_2100_word_offset_0 <= "00000000000000";
    ptr_deref_2287_word_offset_0 <= "00000000000000";
    ptr_deref_2301_word_offset_0 <= "00000000000000";
    type_cast_1193_wire_constant <= "00000000000000000000000000001000";
    type_cast_1218_wire_constant <= "0000000000001000";
    type_cast_1243_wire_constant <= "0000000000001000";
    type_cast_1268_wire_constant <= "0000000000001000";
    type_cast_1293_wire_constant <= "0000000000001000";
    type_cast_1318_wire_constant <= "0000000000001000";
    type_cast_1343_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1368_wire_constant <= "0000000000001000";
    type_cast_1409_wire_constant <= "00000000000000000000000000000011";
    type_cast_1437_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1443_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1472_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1478_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1485_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1496_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1515_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1533_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1551_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1569_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1587_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1605_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1623_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1645_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1664_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1670_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1678_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1690_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1695_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1701_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1714_wire_constant <= "00000000000000000000000000000001";
    type_cast_1720_wire_constant <= "00000000000000000000000000000110";
    type_cast_1729_wire_constant <= "0000000000000000";
    type_cast_1736_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1743_wire_constant <= "0000000000000001";
    type_cast_1749_wire_constant <= "0000000000000001";
    type_cast_1767_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1794_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1800_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1806_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1857_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1865_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1872_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1885_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1891_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1933_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1939_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1946_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1955_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1976_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1994_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2012_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2030_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2048_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2066_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2084_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2106_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2125_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2131_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2139_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2149_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2156_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_2162_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2175_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2185_wire_constant <= "00000000000000000000000000000110";
    type_cast_2196_wire_constant <= "0000000000000000";
    type_cast_2203_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2208_wire_constant <= "0000000000000001";
    type_cast_2214_wire_constant <= "0000000000000001";
    type_cast_2232_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2259_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_2265_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2271_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2303_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2321_wire_constant <= "1111111111111111";
    type_cast_2336_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2354_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2372_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_2385_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_2436_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2454_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2468_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2478_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_2488_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2498_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2508_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2518_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2528_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    phi_stmt_1490: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1493_wire & type_cast_1496_wire_constant;
      req <= phi_stmt_1490_req_0 & phi_stmt_1490_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1490",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1490_ack_0,
          idata => idata,
          odata => indvar425_1490,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1490
    phi_stmt_1684: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1687_wire & type_cast_1690_wire_constant;
      req <= phi_stmt_1684_req_0 & phi_stmt_1684_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1684",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1684_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_1684,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1684
    phi_stmt_1725: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1729_wire_constant & type_cast_1731_wire;
      req <= phi_stmt_1725_req_0 & phi_stmt_1725_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1725",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1725_ack_0,
          idata => idata,
          odata => nx_x022x_xi_1725,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1725
    phi_stmt_1732: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1736_wire_constant & type_cast_1738_wire;
      req <= phi_stmt_1732_req_0 & phi_stmt_1732_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1732",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1732_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_1732,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1732
    phi_stmt_1786: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1789_wire;
      req(0) <= phi_stmt_1786_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1786",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1786_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_1786,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1786
    phi_stmt_1951: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1955_wire_constant & type_cast_1957_wire;
      req <= phi_stmt_1951_req_0 & phi_stmt_1951_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1951",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1951_ack_0,
          idata => idata,
          odata => indvar411_1951,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1951
    phi_stmt_2145: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2149_wire_constant & type_cast_2151_wire;
      req <= phi_stmt_2145_req_0 & phi_stmt_2145_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2145",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2145_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_2145,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2145
    phi_stmt_2190: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2193_wire & type_cast_2196_wire_constant;
      req <= phi_stmt_2190_req_0 & phi_stmt_2190_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2190",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2190_ack_0,
          idata => idata,
          odata => nx_x022x_xi357_2190,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2190
    phi_stmt_2197: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2200_wire & type_cast_2203_wire_constant;
      req <= phi_stmt_2197_req_0 & phi_stmt_2197_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2197",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2197_ack_0,
          idata => idata,
          odata => elementx_x021x_xi358_2197,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2197
    phi_stmt_2251: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_2254_wire;
      req(0) <= phi_stmt_2251_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2251",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2251_ack_0,
          idata => idata,
          odata => shl8x_xi362x_xlcssa_2251,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2251
    phi_stmt_2350: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2354_wire_constant & type_cast_2356_wire;
      req <= phi_stmt_2350_req_0 & phi_stmt_2350_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2350",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2350_ack_0,
          idata => idata,
          odata => indvar_2350,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2350
    -- flow-through select operator MUX_1486_inst
    umax27_1487 <= tmp25_1474 when (tmp26_1480(0) /=  '0') else type_cast_1485_wire_constant;
    -- flow-through select operator MUX_1665_inst
    umax421_1666 <= tmp419_1439 when (tmp420_1445(0) /=  '0') else type_cast_1664_wire_constant;
    -- flow-through select operator MUX_1947_inst
    umax19_1948 <= tmp17_1935 when (tmp18_1941(0) /=  '0') else type_cast_1946_wire_constant;
    -- flow-through select operator MUX_2126_inst
    umax_2127 <= tmp406_1887 when (tmp407_1893(0) /=  '0') else type_cast_2125_wire_constant;
    addr_of_1503_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1503_final_reg_req_0;
      addr_of_1503_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1503_final_reg_req_1;
      addr_of_1503_final_reg_ack_1<= rack(0);
      addr_of_1503_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1503_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1502_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1819_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1819_final_reg_req_0;
      addr_of_1819_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1819_final_reg_req_1;
      addr_of_1819_final_reg_ack_1<= rack(0);
      addr_of_1819_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1819_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1818_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_1820,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1964_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1964_final_reg_req_0;
      addr_of_1964_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1964_final_reg_req_1;
      addr_of_1964_final_reg_ack_1<= rack(0);
      addr_of_1964_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1964_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1963_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1965,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2284_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2284_final_reg_req_0;
      addr_of_2284_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2284_final_reg_req_1;
      addr_of_2284_final_reg_ack_1<= rack(0);
      addr_of_2284_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2284_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2283_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_2285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1188_inst_req_0;
      type_cast_1188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1188_inst_req_1;
      type_cast_1188_inst_ack_1<= rack(0);
      type_cast_1188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_1189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1201_inst_req_0;
      type_cast_1201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1201_inst_req_1;
      type_cast_1201_inst_ack_1<= rack(0);
      type_cast_1201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1213_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1213_inst_req_0;
      type_cast_1213_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1213_inst_req_1;
      type_cast_1213_inst_ack_1<= rack(0);
      type_cast_1213_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1213_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_1214,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1226_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1226_inst_req_0;
      type_cast_1226_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1226_inst_req_1;
      type_cast_1226_inst_ack_1<= rack(0);
      type_cast_1226_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1226_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1227,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1251_inst_req_0;
      type_cast_1251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1251_inst_req_1;
      type_cast_1251_inst_ack_1<= rack(0);
      type_cast_1251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_1248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1263_inst_req_0;
      type_cast_1263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1263_inst_req_1;
      type_cast_1263_inst_ack_1<= rack(0);
      type_cast_1263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_1260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1276_inst_req_0;
      type_cast_1276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1276_inst_req_1;
      type_cast_1276_inst_ack_1<= rack(0);
      type_cast_1276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_1273,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1277,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1288_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1288_inst_req_0;
      type_cast_1288_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1288_inst_req_1;
      type_cast_1288_inst_ack_1<= rack(0);
      type_cast_1288_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1288_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_1285,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1289,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1301_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1301_inst_req_0;
      type_cast_1301_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1301_inst_req_1;
      type_cast_1301_inst_ack_1<= rack(0);
      type_cast_1301_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1301_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_1298,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_1302,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1313_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1313_inst_req_0;
      type_cast_1313_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1313_inst_req_1;
      type_cast_1313_inst_ack_1<= rack(0);
      type_cast_1313_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1313_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_1310,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1314,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1326_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1326_inst_req_0;
      type_cast_1326_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1326_inst_req_1;
      type_cast_1326_inst_ack_1<= rack(0);
      type_cast_1326_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1326_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_1323,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1327,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1338_inst_req_0;
      type_cast_1338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1338_inst_req_1;
      type_cast_1338_inst_ack_1<= rack(0);
      type_cast_1338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_1335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_1339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1351_inst_req_0;
      type_cast_1351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1351_inst_req_1;
      type_cast_1351_inst_ack_1<= rack(0);
      type_cast_1351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_1348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1363_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1363_inst_req_0;
      type_cast_1363_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1363_inst_req_1;
      type_cast_1363_inst_ack_1<= rack(0);
      type_cast_1363_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1363_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_1360,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1376_inst_req_0;
      type_cast_1376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1376_inst_req_1;
      type_cast_1376_inst_ack_1<= rack(0);
      type_cast_1376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_1373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_1377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1385_inst_req_0;
      type_cast_1385_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1385_inst_req_1;
      type_cast_1385_inst_ack_1<= rack(0);
      type_cast_1385_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1385_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_1386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1389_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1389_inst_req_0;
      type_cast_1389_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1389_inst_req_1;
      type_cast_1389_inst_ack_1<= rack(0);
      type_cast_1389_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1389_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_1390,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1404_inst_req_0;
      type_cast_1404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1404_inst_req_1;
      type_cast_1404_inst_ack_1<= rack(0);
      type_cast_1404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1404_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1403_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_1405,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1432_inst_req_0;
      type_cast_1432_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1432_inst_req_1;
      type_cast_1432_inst_ack_1<= rack(0);
      type_cast_1432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1431_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp418_1433,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1448_inst_req_0;
      type_cast_1448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1448_inst_req_1;
      type_cast_1448_inst_ack_1<= rack(0);
      type_cast_1448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1449,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1457_inst_req_0;
      type_cast_1457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1457_inst_req_1;
      type_cast_1457_inst_ack_1<= rack(0);
      type_cast_1457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp22_1458,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1467_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1467_inst_req_0;
      type_cast_1467_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1467_inst_req_1;
      type_cast_1467_inst_ack_1<= rack(0);
      type_cast_1467_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1467_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1466_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_1468,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1493_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1493_inst_req_0;
      type_cast_1493_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1493_inst_req_1;
      type_cast_1493_inst_ack_1<= rack(0);
      type_cast_1493_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1493_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext426_1647,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1493_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1510_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1510_inst_req_0;
      type_cast_1510_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1510_inst_req_1;
      type_cast_1510_inst_ack_1<= rack(0);
      type_cast_1510_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1510_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_1507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1511,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1523_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1523_inst_req_0;
      type_cast_1523_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1523_inst_req_1;
      type_cast_1523_inst_ack_1<= rack(0);
      type_cast_1523_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1523_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_1520,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_1524,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1541_inst_req_0;
      type_cast_1541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1541_inst_req_1;
      type_cast_1541_inst_ack_1<= rack(0);
      type_cast_1541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_1538,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_1542,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1559_inst_req_0;
      type_cast_1559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1559_inst_req_1;
      type_cast_1559_inst_ack_1<= rack(0);
      type_cast_1559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_1556,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1560,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1577_inst_req_0;
      type_cast_1577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1577_inst_req_1;
      type_cast_1577_inst_ack_1<= rack(0);
      type_cast_1577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_1574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_1578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1595_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1595_inst_req_0;
      type_cast_1595_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1595_inst_req_1;
      type_cast_1595_inst_ack_1<= rack(0);
      type_cast_1595_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1595_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_1592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_1596,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1613_inst_req_0;
      type_cast_1613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1613_inst_req_1;
      type_cast_1613_inst_ack_1<= rack(0);
      type_cast_1613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_1610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_1614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1631_inst_req_0;
      type_cast_1631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1631_inst_req_1;
      type_cast_1631_inst_ack_1<= rack(0);
      type_cast_1631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_1628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_1632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1675_inst
    process(tmp422_1672) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp422_1672(63 downto 0);
      type_cast_1675_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1680_inst
    process(ASHR_i64_i64_1679_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1679_wire(63 downto 0);
      phitmp_1681 <= tmp_var; -- 
    end process;
    type_cast_1687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1687_inst_req_0;
      type_cast_1687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1687_inst_req_1;
      type_cast_1687_inst_ack_1<= rack(0);
      type_cast_1687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_1681,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1687_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1731_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1731_inst_req_0;
      type_cast_1731_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1731_inst_req_1;
      type_cast_1731_inst_ack_1<= rack(0);
      type_cast_1731_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1731_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_35_1751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1731_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1738_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1738_inst_req_0;
      type_cast_1738_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1738_inst_req_1;
      type_cast_1738_inst_ack_1<= rack(0);
      type_cast_1738_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1738_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1738_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1757_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1757_inst_req_0;
      type_cast_1757_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1757_inst_req_1;
      type_cast_1757_inst_ack_1<= rack(0);
      type_cast_1757_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1757_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1754,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1758,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1772_inst_req_0;
      type_cast_1772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1772_inst_req_1;
      type_cast_1772_inst_ack_1<= rack(0);
      type_cast_1772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1745,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1789_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1789_inst_req_0;
      type_cast_1789_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1789_inst_req_1;
      type_cast_1789_inst_ack_1<= rack(0);
      type_cast_1789_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1789_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1789_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1829_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1829_inst_req_0;
      type_cast_1829_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1829_inst_req_1;
      type_cast_1829_inst_ack_1<= rack(0);
      type_cast_1829_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1829_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1830,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1833_inst_req_0;
      type_cast_1833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1833_inst_req_1;
      type_cast_1833_inst_ack_1<= rack(0);
      type_cast_1833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_1382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_1834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1837_inst_req_0;
      type_cast_1837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1837_inst_req_1;
      type_cast_1837_inst_ack_1<= rack(0);
      type_cast_1837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1837_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1838,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1862_inst
    process(sext_1859) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1859(63 downto 0);
      type_cast_1862_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1867_inst
    process(ASHR_i64_i64_1866_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1866_wire(63 downto 0);
      conv155_1868 <= tmp_var; -- 
    end process;
    type_cast_1896_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1896_inst_req_0;
      type_cast_1896_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1896_inst_req_1;
      type_cast_1896_inst_ack_1<= rack(0);
      type_cast_1896_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1896_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp9_1897,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1905_inst_req_0;
      type_cast_1905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1905_inst_req_1;
      type_cast_1905_inst_ack_1<= rack(0);
      type_cast_1905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp11_1906,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1914_inst_req_0;
      type_cast_1914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1914_inst_req_1;
      type_cast_1914_inst_ack_1<= rack(0);
      type_cast_1914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_1382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1923_inst_req_0;
      type_cast_1923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1923_inst_req_1;
      type_cast_1923_inst_ack_1<= rack(0);
      type_cast_1923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_1920,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_1924,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1928_inst_req_0;
      type_cast_1928_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1928_inst_req_1;
      type_cast_1928_inst_ack_1<= rack(0);
      type_cast_1928_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1927_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp16_1929,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1957_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1957_inst_req_0;
      type_cast_1957_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1957_inst_req_1;
      type_cast_1957_inst_ack_1<= rack(0);
      type_cast_1957_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1957_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext412_2108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1957_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1971_inst_req_0;
      type_cast_1971_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1971_inst_req_1;
      type_cast_1971_inst_ack_1<= rack(0);
      type_cast_1971_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1971_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_1968,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1972,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1984_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1984_inst_req_0;
      type_cast_1984_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1984_inst_req_1;
      type_cast_1984_inst_ack_1<= rack(0);
      type_cast_1984_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1984_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1981,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1985,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2002_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2002_inst_req_0;
      type_cast_2002_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2002_inst_req_1;
      type_cast_2002_inst_ack_1<= rack(0);
      type_cast_2002_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2002_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1999,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_2003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2020_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2020_inst_req_0;
      type_cast_2020_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2020_inst_req_1;
      type_cast_2020_inst_ack_1<= rack(0);
      type_cast_2020_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2020_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_2017,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_2021,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2038_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2038_inst_req_0;
      type_cast_2038_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2038_inst_req_1;
      type_cast_2038_inst_ack_1<= rack(0);
      type_cast_2038_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2038_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_2035,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_2039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2056_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2056_inst_req_0;
      type_cast_2056_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2056_inst_req_1;
      type_cast_2056_inst_ack_1<= rack(0);
      type_cast_2056_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2056_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_2053,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_2057,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2074_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2074_inst_req_0;
      type_cast_2074_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2074_inst_req_1;
      type_cast_2074_inst_ack_1<= rack(0);
      type_cast_2074_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2074_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_2071,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_2075,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2092_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2092_inst_req_0;
      type_cast_2092_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2092_inst_req_1;
      type_cast_2092_inst_ack_1<= rack(0);
      type_cast_2092_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2092_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_2089,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_2093,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2136_inst
    process(tmp408_2133) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp408_2133(63 downto 0);
      type_cast_2136_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2141_inst
    process(ASHR_i64_i64_2140_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_2140_wire(63 downto 0);
      phitmp387_2142 <= tmp_var; -- 
    end process;
    type_cast_2151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2151_inst_req_0;
      type_cast_2151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2151_inst_req_1;
      type_cast_2151_inst_ack_1<= rack(0);
      type_cast_2151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp387_2142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2151_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2180_inst_req_0;
      type_cast_2180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2180_inst_req_1;
      type_cast_2180_inst_ack_1<= rack(0);
      type_cast_2180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_59_2177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi354_2181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2193_inst_req_0;
      type_cast_2193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2193_inst_req_1;
      type_cast_2193_inst_ack_1<= rack(0);
      type_cast_2193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_71_2216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2193_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2200_inst_req_0;
      type_cast_2200_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2200_inst_req_1;
      type_cast_2200_inst_ack_1<= rack(0);
      type_cast_2200_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2200_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi362_2234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2200_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2222_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2222_inst_req_0;
      type_cast_2222_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2222_inst_req_1;
      type_cast_2222_inst_ack_1<= rack(0);
      type_cast_2222_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2222_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi359_2219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi360_2223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2237_inst_req_0;
      type_cast_2237_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2237_inst_req_1;
      type_cast_2237_inst_ack_1<= rack(0);
      type_cast_2237_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2237_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp388_2210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi363_2238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2254_inst_req_0;
      type_cast_2254_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2254_inst_req_1;
      type_cast_2254_inst_ack_1<= rack(0);
      type_cast_2254_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2254_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi362_2234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2254_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2331_inst_req_0;
      type_cast_2331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2331_inst_req_1;
      type_cast_2331_inst_ack_1<= rack(0);
      type_cast_2331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp389_2323,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_2332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2341_inst_req_0;
      type_cast_2341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2341_inst_req_1;
      type_cast_2341_inst_ack_1<= rack(0);
      type_cast_2341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp393_2328,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_2342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2356_inst_req_0;
      type_cast_2356_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2356_inst_req_1;
      type_cast_2356_inst_ack_1<= rack(0);
      type_cast_2356_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2387,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2356_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2403_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2403_inst_req_0;
      type_cast_2403_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2403_inst_req_1;
      type_cast_2403_inst_ack_1<= rack(0);
      type_cast_2403_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2403_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2402_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_2404,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2418_inst_req_0;
      type_cast_2418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2418_inst_req_1;
      type_cast_2418_inst_ack_1<= rack(0);
      type_cast_2418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2417_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_2419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2427_inst_req_0;
      type_cast_2427_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2427_inst_req_1;
      type_cast_2427_inst_ack_1<= rack(0);
      type_cast_2427_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2427_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add43_1307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv281_2428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2431_inst_req_0;
      type_cast_2431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2431_inst_req_1;
      type_cast_2431_inst_ack_1<= rack(0);
      type_cast_2431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_1282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv283_2432,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2451_inst
    process(sext352_2448) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext352_2448(63 downto 0);
      type_cast_2451_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2456_inst
    process(ASHR_i64_i64_2455_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_2455_wire(63 downto 0);
      conv288_2457 <= tmp_var; -- 
    end process;
    type_cast_2463_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2463_inst_req_0;
      type_cast_2463_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2463_inst_req_1;
      type_cast_2463_inst_ack_1<= rack(0);
      type_cast_2463_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2463_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_2424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv292_2464,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2473_inst_req_0;
      type_cast_2473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2473_inst_req_1;
      type_cast_2473_inst_ack_1<= rack(0);
      type_cast_2473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr295_2470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv298_2474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2483_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2483_inst_req_0;
      type_cast_2483_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2483_inst_req_1;
      type_cast_2483_inst_ack_1<= rack(0);
      type_cast_2483_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2483_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr301_2480,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv304_2484,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2493_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2493_inst_req_0;
      type_cast_2493_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2493_inst_req_1;
      type_cast_2493_inst_ack_1<= rack(0);
      type_cast_2493_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2493_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr307_2490,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv310_2494,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2503_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2503_inst_req_0;
      type_cast_2503_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2503_inst_req_1;
      type_cast_2503_inst_ack_1<= rack(0);
      type_cast_2503_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2503_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr313_2500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv316_2504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2513_inst_req_0;
      type_cast_2513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2513_inst_req_1;
      type_cast_2513_inst_ack_1<= rack(0);
      type_cast_2513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr319_2510,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_2514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2523_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2523_inst_req_0;
      type_cast_2523_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2523_inst_req_1;
      type_cast_2523_inst_ack_1<= rack(0);
      type_cast_2523_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2523_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr325_2520,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv328_2524,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2533_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2533_inst_req_0;
      type_cast_2533_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2533_inst_req_1;
      type_cast_2533_inst_ack_1<= rack(0);
      type_cast_2533_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2533_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr331_2530,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv334_2534,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1502_index_1_rename
    process(R_indvar425_1501_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar425_1501_resized;
      ov(13 downto 0) := iv;
      R_indvar425_1501_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1502_index_1_resize
    process(indvar425_1490) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar425_1490;
      ov := iv(13 downto 0);
      R_indvar425_1501_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1502_root_address_inst
    process(array_obj_ref_1502_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1502_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1502_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1818_index_1_rename
    process(R_ix_x0x_xlcssa_1817_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1817_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1817_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1818_index_1_resize
    process(ix_x0x_xlcssa_1684) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_1684;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1817_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1818_root_address_inst
    process(array_obj_ref_1818_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1818_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1818_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1963_index_1_rename
    process(R_indvar411_1962_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar411_1962_resized;
      ov(13 downto 0) := iv;
      R_indvar411_1962_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1963_index_1_resize
    process(indvar411_1951) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar411_1951;
      ov := iv(13 downto 0);
      R_indvar411_1962_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1963_root_address_inst
    process(array_obj_ref_1963_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1963_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1963_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2283_index_1_rename
    process(R_ix_x1x_xlcssa_2282_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_2282_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_2282_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2283_index_1_resize
    process(ix_x1x_xlcssa_2145) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_2145;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_2282_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2283_root_address_inst
    process(array_obj_ref_2283_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2283_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2283_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1639_addr_0
    process(ptr_deref_1639_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1639_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1639_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1639_base_resize
    process(arrayidx_1504) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1504;
      ov := iv(13 downto 0);
      ptr_deref_1639_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1639_gather_scatter
    process(add132_1637) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_1637;
      ov(63 downto 0) := iv;
      ptr_deref_1639_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1639_root_address_inst
    process(ptr_deref_1639_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1639_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1639_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1822_addr_0
    process(ptr_deref_1822_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1822_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1822_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1822_base_resize
    process(arrayidx143_1820) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_1820;
      ov := iv(13 downto 0);
      ptr_deref_1822_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1822_gather_scatter
    process(shl14x_xi_1813) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_1813;
      ov(63 downto 0) := iv;
      ptr_deref_1822_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1822_root_address_inst
    process(ptr_deref_1822_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1822_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1822_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_addr_0
    process(ptr_deref_2100_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2100_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2100_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_base_resize
    process(arrayidx211_1965) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1965;
      ov := iv(13 downto 0);
      ptr_deref_2100_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_gather_scatter
    process(add207_2098) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_2098;
      ov(63 downto 0) := iv;
      ptr_deref_2100_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_root_address_inst
    process(ptr_deref_2100_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2100_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2100_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2287_addr_0
    process(ptr_deref_2287_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2287_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2287_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2287_base_resize
    process(arrayidx226_2285) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_2285;
      ov := iv(13 downto 0);
      ptr_deref_2287_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2287_gather_scatter
    process(shl14x_xi372_2278) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi372_2278;
      ov(63 downto 0) := iv;
      ptr_deref_2287_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2287_root_address_inst
    process(ptr_deref_2287_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2287_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2287_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2301_addr_0
    process(ptr_deref_2301_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2301_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2301_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2301_base_resize
    process(iNsTr_48_2299) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_48_2299;
      ov := iv(13 downto 0);
      ptr_deref_2301_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2301_gather_scatter
    process(type_cast_2303_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_2303_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_2301_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2301_root_address_inst
    process(ptr_deref_2301_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2301_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2301_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1412_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp383_1411;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1412_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1412_branch_req_0,
          ack0 => if_stmt_1412_branch_ack_0,
          ack1 => if_stmt_1412_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1653_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond28_1652;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1653_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1653_branch_req_0,
          ack0 => if_stmt_1653_branch_ack_0,
          ack1 => if_stmt_1653_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1704_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1703;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1704_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1704_branch_req_0,
          ack0 => if_stmt_1704_branch_ack_0,
          ack1 => if_stmt_1704_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1779_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1778;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1779_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1779_branch_req_0,
          ack0 => if_stmt_1779_branch_ack_0,
          ack1 => if_stmt_1779_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1875_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161379_1874;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1875_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1875_branch_req_0,
          ack0 => if_stmt_1875_branch_ack_0,
          ack1 => if_stmt_1875_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2114_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_2113;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2114_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2114_branch_req_0,
          ack0 => if_stmt_2114_branch_ack_0,
          ack1 => if_stmt_2114_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2165_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_2164;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2165_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2165_branch_req_0,
          ack0 => if_stmt_2165_branch_ack_0,
          ack1 => if_stmt_2165_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2244_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi364_2243;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2244_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2244_branch_req_0,
          ack0 => if_stmt_2244_branch_ack_0,
          ack1 => if_stmt_2244_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2393_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_2392;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2393_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2393_branch_req_0,
          ack0 => if_stmt_2393_branch_ack_0,
          ack1 => if_stmt_2393_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1744_inst
    process(nx_x022x_xi_1725) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_1725, type_cast_1743_wire_constant, tmp_var);
      tmp_1745 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1750_inst
    process(nx_x022x_xi_1725) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_1725, type_cast_1749_wire_constant, tmp_var);
      iNsTr_35_1751 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2209_inst
    process(nx_x022x_xi357_2190) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi357_2190, type_cast_2208_wire_constant, tmp_var);
      tmp388_2210 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2215_inst
    process(nx_x022x_xi357_2190) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi357_2190, type_cast_2214_wire_constant, tmp_var);
      iNsTr_71_2216 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2322_inst
    process(add53_1332) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_1332, type_cast_2321_wire_constant, tmp_var);
      tmp389_2323 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1646_inst
    process(indvar425_1490) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar425_1490, type_cast_1645_wire_constant, tmp_var);
      indvarx_xnext426_1647 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2107_inst
    process(indvar411_1951) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar411_1951, type_cast_2106_wire_constant, tmp_var);
      indvarx_xnext412_2108 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2337_inst
    process(tmp3_2332) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_2332, type_cast_2336_wire_constant, tmp_var);
      tmp4_2338 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2386_inst
    process(indvar_2350) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2350, type_cast_2385_wire_constant, tmp_var);
      indvarx_xnext_2387 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1721_inst
    process(conv2x_xi_1716) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_1716, type_cast_1720_wire_constant, tmp_var);
      shlx_xi_1722 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2186_inst
    process(conv2x_xi354_2181) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi354_2181, type_cast_2185_wire_constant, tmp_var);
      shlx_xi355_2187 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1696_inst
    process(conv83_1405) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_1405, type_cast_1695_wire_constant, tmp_var);
      and_1697 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1801_inst
    process(Bx_xnot_1796) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1796, type_cast_1800_wire_constant, tmp_var);
      add1216x_xi_1802 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2157_inst
    process(conv155_1868) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_1868, type_cast_2156_wire_constant, tmp_var);
      and217_2158 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2266_inst
    process(iNsTr_97_2261) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_97_2261, type_cast_2265_wire_constant, tmp_var);
      add1216x_xi370_2267 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2373_inst
    process(mul253_2362) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul253_2362, type_cast_2372_wire_constant, tmp_var);
      conv254_2374 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1679_inst
    process(type_cast_1675_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1675_wire, type_cast_1678_wire_constant, tmp_var);
      ASHR_i64_i64_1679_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1866_inst
    process(type_cast_1862_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1862_wire, type_cast_1865_wire_constant, tmp_var);
      ASHR_i64_i64_1866_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_2140_inst
    process(type_cast_2136_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2136_wire, type_cast_2139_wire_constant, tmp_var);
      ASHR_i64_i64_2140_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_2455_inst
    process(type_cast_2451_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2451_wire, type_cast_2454_wire_constant, tmp_var);
      ASHR_i64_i64_2455_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1651_inst
    process(indvarx_xnext426_1647, umax27_1487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext426_1647, umax27_1487, tmp_var);
      exitcond28_1652 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1702_inst
    process(and_1697) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_1697, type_cast_1701_wire_constant, tmp_var);
      tobool_1703 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2112_inst
    process(indvarx_xnext412_2108, umax19_1948) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext412_2108, umax19_1948, tmp_var);
      exitcond_2113 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2163_inst
    process(and217_2158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_2158, type_cast_2162_wire_constant, tmp_var);
      tobool218_2164 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_2391_inst
    process(indvarx_xnext_2387, tmp4_2338) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_2387, tmp4_2338, tmp_var);
      exitcond5_2392 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1438_inst
    process(tmp418_1433) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp418_1433, type_cast_1437_wire_constant, tmp_var);
      tmp419_1439 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1473_inst
    process(tmp24_1468) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp24_1468, type_cast_1472_wire_constant, tmp_var);
      tmp25_1474 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1886_inst
    process(conv155_1868) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1868, type_cast_1885_wire_constant, tmp_var);
      tmp406_1887 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1934_inst
    process(tmp16_1929) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp16_1929, type_cast_1933_wire_constant, tmp_var);
      tmp17_1935 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2469_inst
    process(sub_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2424, type_cast_2468_wire_constant, tmp_var);
      shr295_2470 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2479_inst
    process(sub_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2424, type_cast_2478_wire_constant, tmp_var);
      shr301_2480 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2489_inst
    process(sub_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2424, type_cast_2488_wire_constant, tmp_var);
      shr307_2490 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2499_inst
    process(sub_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2424, type_cast_2498_wire_constant, tmp_var);
      shr313_2500 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2509_inst
    process(sub_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2424, type_cast_2508_wire_constant, tmp_var);
      shr319_2510 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2519_inst
    process(sub_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2424, type_cast_2518_wire_constant, tmp_var);
      shr325_2520 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2529_inst
    process(sub_2424) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_2424, type_cast_2528_wire_constant, tmp_var);
      shr331_2530 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2327_inst
    process(add73_1382, add23_1257) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1382, add23_1257, tmp_var);
      tmp393_2328 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1394_inst
    process(conv79_1386, add_1207) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_1386, add_1207, tmp_var);
      mul_1395 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1399_inst
    process(mul_1395, conv81_1390) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1395, conv81_1390, tmp_var);
      mul82_1400 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1422_inst
    process(add_1207, conv79_1386) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1207, conv79_1386, tmp_var);
      tmp415_1423 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1427_inst
    process(tmp415_1423, conv81_1390) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp415_1423, conv81_1390, tmp_var);
      tmp417_1428 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1453_inst
    process(add_1207, tmp20_1449) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1207, tmp20_1449, tmp_var);
      tmp21_1454 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1462_inst
    process(tmp21_1454, tmp22_1458) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp21_1454, tmp22_1458, tmp_var);
      tmp23_1463 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1842_inst
    process(conv153_1838, conv145_1830) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_1838, conv145_1830, tmp_var);
      mul148_1843 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1847_inst
    process(mul148_1843, add63_1357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_1843, add63_1357, tmp_var);
      mul151_1848 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1852_inst
    process(mul151_1848, conv147_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_1848, conv147_1834, tmp_var);
      mul154_1853 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1901_inst
    process(add63_1357, tmp9_1897) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_1357, tmp9_1897, tmp_var);
      tmp10_1902 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1910_inst
    process(tmp10_1902, tmp11_1906) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp10_1902, tmp11_1906, tmp_var);
      tmp12_1911 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1919_inst
    process(tmp12_1911, tmp13_1915) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_1911, tmp13_1915, tmp_var);
      tmp14_1920 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2346_inst
    process(add63_1357, tmp6_2342) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_1357, tmp6_2342, tmp_var);
      tmp7_2347 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2361_inst
    process(tmp7_2347, indvar_2350) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp7_2347, indvar_2350, tmp_var);
      mul253_2362 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2442_inst
    process(mul284_2438, conv281_2428) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul284_2438, conv281_2428, tmp_var);
      mul287_2443 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2447_inst
    process(mul287_2443, conv153_1838) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul287_2443, conv153_1838, tmp_var);
      sext352_2448 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1231_inst
    process(shl10_1220, conv12_1227) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_1220, conv12_1227, tmp_var);
      add13_1232 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1256_inst
    process(shl20_1245, conv22_1252) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_1245, conv22_1252, tmp_var);
      add23_1257 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1281_inst
    process(shl30_1270, conv32_1277) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_1270, conv32_1277, tmp_var);
      add33_1282 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1306_inst
    process(shl40_1295, conv42_1302) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_1295, conv42_1302, tmp_var);
      add43_1307 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1331_inst
    process(shl50_1320, conv52_1327) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_1320, conv52_1327, tmp_var);
      add53_1332 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1381_inst
    process(shl70_1370, conv72_1377) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_1370, conv72_1377, tmp_var);
      add73_1382 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1206_inst
    process(shl_1195, conv3_1202) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1195, conv3_1202, tmp_var);
      add_1207 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1356_inst
    process(shl60_1345, conv62_1352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_1345, conv62_1352, tmp_var);
      add63_1357 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1528_inst
    process(shl92_1517, conv95_1524) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_1517, conv95_1524, tmp_var);
      add96_1529 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1546_inst
    process(shl98_1535, conv101_1542) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_1535, conv101_1542, tmp_var);
      add102_1547 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1564_inst
    process(shl104_1553, conv107_1560) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_1553, conv107_1560, tmp_var);
      add108_1565 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1582_inst
    process(shl110_1571, conv113_1578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_1571, conv113_1578, tmp_var);
      add114_1583 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1600_inst
    process(shl116_1589, conv119_1596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_1589, conv119_1596, tmp_var);
      add120_1601 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1618_inst
    process(shl122_1607, conv125_1614) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_1607, conv125_1614, tmp_var);
      add126_1619 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1636_inst
    process(shl128_1625, conv131_1632) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_1625, conv131_1632, tmp_var);
      add132_1637 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1762_inst
    process(conv5x_xi_1758, elementx_x021x_xi_1732) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1758, elementx_x021x_xi_1732, tmp_var);
      addx_xi_1763 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1989_inst
    process(shl167_1978, conv170_1985) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1978, conv170_1985, tmp_var);
      add171_1990 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2007_inst
    process(shl173_1996, conv176_2003) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1996, conv176_2003, tmp_var);
      add177_2008 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2025_inst
    process(shl179_2014, conv182_2021) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_2014, conv182_2021, tmp_var);
      add183_2026 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2043_inst
    process(shl185_2032, conv188_2039) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_2032, conv188_2039, tmp_var);
      add189_2044 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2061_inst
    process(shl191_2050, conv194_2057) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_2050, conv194_2057, tmp_var);
      add195_2062 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2079_inst
    process(shl197_2068, conv200_2075) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_2068, conv200_2075, tmp_var);
      add201_2080 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2097_inst
    process(shl203_2086, conv206_2093) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_2086, conv206_2093, tmp_var);
      add207_2098 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2227_inst
    process(conv5x_xi360_2223, elementx_x021x_xi358_2197) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi360_2223, elementx_x021x_xi358_2197, tmp_var);
      addx_xi361_2228 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1219_inst
    process(conv9_1214) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_1214, type_cast_1218_wire_constant, tmp_var);
      shl10_1220 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1244_inst
    process(conv19_1239) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_1239, type_cast_1243_wire_constant, tmp_var);
      shl20_1245 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1269_inst
    process(conv29_1264) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_1264, type_cast_1268_wire_constant, tmp_var);
      shl30_1270 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1294_inst
    process(conv39_1289) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_1289, type_cast_1293_wire_constant, tmp_var);
      shl40_1295 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1319_inst
    process(conv49_1314) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1314, type_cast_1318_wire_constant, tmp_var);
      shl50_1320 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1369_inst
    process(conv69_1364) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_1364, type_cast_1368_wire_constant, tmp_var);
      shl70_1370 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1194_inst
    process(conv1_1189) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_1189, type_cast_1193_wire_constant, tmp_var);
      shl_1195 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1715_inst
    process(mul82_1400) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_1400, type_cast_1714_wire_constant, tmp_var);
      conv2x_xi_1716 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1344_inst
    process(conv59_1339) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_1339, type_cast_1343_wire_constant, tmp_var);
      shl60_1345 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1516_inst
    process(conv90_1511) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_1511, type_cast_1515_wire_constant, tmp_var);
      shl92_1517 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1534_inst
    process(add96_1529) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_1529, type_cast_1533_wire_constant, tmp_var);
      shl98_1535 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1552_inst
    process(add102_1547) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_1547, type_cast_1551_wire_constant, tmp_var);
      shl104_1553 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1570_inst
    process(add108_1565) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_1565, type_cast_1569_wire_constant, tmp_var);
      shl110_1571 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1588_inst
    process(add114_1583) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_1583, type_cast_1587_wire_constant, tmp_var);
      shl116_1589 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1606_inst
    process(add120_1601) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_1601, type_cast_1605_wire_constant, tmp_var);
      shl122_1607 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1624_inst
    process(add126_1619) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_1619, type_cast_1623_wire_constant, tmp_var);
      shl128_1625 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1671_inst
    process(umax421_1666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax421_1666, type_cast_1670_wire_constant, tmp_var);
      tmp422_1672 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1768_inst
    process(addx_xi_1763) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1763, type_cast_1767_wire_constant, tmp_var);
      shl8x_xi_1769 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1795_inst
    process(conv83_1405) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_1405, type_cast_1794_wire_constant, tmp_var);
      Bx_xnot_1796 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1812_inst
    process(shl8x_xix_xlcssa_1786, sh_promx_xi_1808) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_1786, sh_promx_xi_1808, tmp_var);
      shl14x_xi_1813 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1858_inst
    process(mul154_1853) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1853, type_cast_1857_wire_constant, tmp_var);
      sext_1859 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1977_inst
    process(conv165_1972) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_1972, type_cast_1976_wire_constant, tmp_var);
      shl167_1978 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1995_inst
    process(add171_1990) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1990, type_cast_1994_wire_constant, tmp_var);
      shl173_1996 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2013_inst
    process(add177_2008) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_2008, type_cast_2012_wire_constant, tmp_var);
      shl179_2014 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2031_inst
    process(add183_2026) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_2026, type_cast_2030_wire_constant, tmp_var);
      shl185_2032 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2049_inst
    process(add189_2044) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_2044, type_cast_2048_wire_constant, tmp_var);
      shl191_2050 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2067_inst
    process(add195_2062) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_2062, type_cast_2066_wire_constant, tmp_var);
      shl197_2068 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2085_inst
    process(add201_2080) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_2080, type_cast_2084_wire_constant, tmp_var);
      shl203_2086 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2132_inst
    process(umax_2127) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_2127, type_cast_2131_wire_constant, tmp_var);
      tmp408_2133 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2176_inst
    process(mul154_1853) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1853, type_cast_2175_wire_constant, tmp_var);
      iNsTr_59_2177 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2233_inst
    process(addx_xi361_2228) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi361_2228, type_cast_2232_wire_constant, tmp_var);
      shl8x_xi362_2234 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2260_inst
    process(mul154_1853) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1853, type_cast_2259_wire_constant, tmp_var);
      iNsTr_97_2261 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2277_inst
    process(shl8x_xi362x_xlcssa_2251, sh_promx_xi371_2273) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi362x_xlcssa_2251, sh_promx_xi371_2273, tmp_var);
      shl14x_xi372_2278 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_2437_inst
    process(conv283_2432) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv283_2432, type_cast_2436_wire_constant, tmp_var);
      mul284_2438 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_2423_inst
    process(conv276_2419, conv230_2404) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv276_2419, conv230_2404, tmp_var);
      sub_2424 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1410_inst
    process(mul82_1400) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_1400, type_cast_1409_wire_constant, tmp_var);
      cmp383_1411 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1444_inst
    process(tmp419_1439) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp419_1439, type_cast_1443_wire_constant, tmp_var);
      tmp420_1445 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1479_inst
    process(tmp25_1474) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp25_1474, type_cast_1478_wire_constant, tmp_var);
      tmp26_1480 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1873_inst
    process(conv155_1868) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_1868, type_cast_1872_wire_constant, tmp_var);
      cmp161379_1874 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1892_inst
    process(tmp406_1887) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp406_1887, type_cast_1891_wire_constant, tmp_var);
      tmp407_1893 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1940_inst
    process(tmp17_1935) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp17_1935, type_cast_1939_wire_constant, tmp_var);
      tmp18_1941 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1777_inst
    process(convx_xi_1773, shlx_xi_1722) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1773, shlx_xi_1722, tmp_var);
      cmpx_xi_1778 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2242_inst
    process(convx_xi363_2238, shlx_xi355_2187) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi363_2238, shlx_xi355_2187, tmp_var);
      cmpx_xi364_2243 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1807_inst
    process(add1216x_xi_1802) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_1802, type_cast_1806_wire_constant, tmp_var);
      sh_promx_xi_1808 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_2272_inst
    process(add1216x_xi370_2267) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi370_2267, type_cast_2271_wire_constant, tmp_var);
      sh_promx_xi371_2273 <= tmp_var; --
    end process;
    -- shared split operator group (122) : array_obj_ref_1502_index_offset 
    ApIntAdd_group_122: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar425_1501_scaled;
      array_obj_ref_1502_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1502_index_offset_req_0;
      array_obj_ref_1502_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1502_index_offset_req_1;
      array_obj_ref_1502_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_122_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_122_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- shared split operator group (123) : array_obj_ref_1818_index_offset 
    ApIntAdd_group_123: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1817_scaled;
      array_obj_ref_1818_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1818_index_offset_req_0;
      array_obj_ref_1818_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1818_index_offset_req_1;
      array_obj_ref_1818_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_123_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_123_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : array_obj_ref_1963_index_offset 
    ApIntAdd_group_124: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar411_1962_scaled;
      array_obj_ref_1963_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1963_index_offset_req_0;
      array_obj_ref_1963_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1963_index_offset_req_1;
      array_obj_ref_1963_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_124_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_124_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : array_obj_ref_2283_index_offset 
    ApIntAdd_group_125: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_2282_scaled;
      array_obj_ref_2283_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2283_index_offset_req_0;
      array_obj_ref_2283_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2283_index_offset_req_1;
      array_obj_ref_2283_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_125_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_125_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- unary operator type_cast_1403_inst
    process(mul82_1400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_1400, tmp_var);
      type_cast_1403_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1431_inst
    process(tmp417_1428) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp417_1428, tmp_var);
      type_cast_1431_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1466_inst
    process(tmp23_1463) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp23_1463, tmp_var);
      type_cast_1466_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1927_inst
    process(tmp15_1924) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp15_1924, tmp_var);
      type_cast_1927_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2402_inst
    process(call229_2307) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_2307, tmp_var);
      type_cast_2402_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2417_inst
    process(call275_2414) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_2414, tmp_var);
      type_cast_2417_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1639_store_0 ptr_deref_1822_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1639_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1822_store_0_req_0;
      ptr_deref_1639_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1822_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1639_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1822_store_0_req_1;
      ptr_deref_1639_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1822_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1639_word_address_0 & ptr_deref_1822_word_address_0;
      data_in <= ptr_deref_1639_data_0 & ptr_deref_1822_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 4,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_2100_store_0 ptr_deref_2287_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2100_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2287_store_0_req_0;
      ptr_deref_2100_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2287_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2100_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2287_store_0_req_1;
      ptr_deref_2100_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2287_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2100_word_address_0 & ptr_deref_2287_word_address_0;
      data_in <= ptr_deref_2100_data_0 & ptr_deref_2287_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_2301_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2301_store_0_req_0;
      ptr_deref_2301_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2301_store_0_req_1;
      ptr_deref_2301_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2301_word_address_0;
      data_in <= ptr_deref_2301_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_input_done_pipe_2406_inst RPIPE_input_done_pipe_2410_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_input_done_pipe_2406_inst_req_0;
      reqL_unguarded(0) <= RPIPE_input_done_pipe_2410_inst_req_0;
      RPIPE_input_done_pipe_2406_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_input_done_pipe_2410_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_input_done_pipe_2406_inst_req_1;
      reqR_unguarded(0) <= RPIPE_input_done_pipe_2410_inst_req_1;
      RPIPE_input_done_pipe_2406_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_input_done_pipe_2410_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      call270_2407 <= data_out(15 downto 8);
      call273_2411 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_maxpool_input_pipe_1555_inst RPIPE_maxpool_input_pipe_1506_inst RPIPE_maxpool_input_pipe_1967_inst RPIPE_maxpool_input_pipe_2016_inst RPIPE_maxpool_input_pipe_1998_inst RPIPE_maxpool_input_pipe_2070_inst RPIPE_maxpool_input_pipe_1519_inst RPIPE_maxpool_input_pipe_1573_inst RPIPE_maxpool_input_pipe_1627_inst RPIPE_maxpool_input_pipe_1537_inst RPIPE_maxpool_input_pipe_1591_inst RPIPE_maxpool_input_pipe_2088_inst RPIPE_maxpool_input_pipe_1980_inst RPIPE_maxpool_input_pipe_1753_inst RPIPE_maxpool_input_pipe_1609_inst RPIPE_maxpool_input_pipe_2218_inst RPIPE_maxpool_input_pipe_2034_inst RPIPE_maxpool_input_pipe_1184_inst RPIPE_maxpool_input_pipe_1197_inst RPIPE_maxpool_input_pipe_1209_inst RPIPE_maxpool_input_pipe_1222_inst RPIPE_maxpool_input_pipe_1234_inst RPIPE_maxpool_input_pipe_1247_inst RPIPE_maxpool_input_pipe_1259_inst RPIPE_maxpool_input_pipe_1272_inst RPIPE_maxpool_input_pipe_1284_inst RPIPE_maxpool_input_pipe_2052_inst RPIPE_maxpool_input_pipe_1297_inst RPIPE_maxpool_input_pipe_1309_inst RPIPE_maxpool_input_pipe_1322_inst RPIPE_maxpool_input_pipe_1334_inst RPIPE_maxpool_input_pipe_1347_inst RPIPE_maxpool_input_pipe_1359_inst RPIPE_maxpool_input_pipe_1372_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_1555_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_1506_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_1967_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_2016_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_1998_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_2070_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_1519_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_1573_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_1627_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_1537_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_1591_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_2088_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_1980_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_1753_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_1609_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_2218_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_2034_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_1184_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_1197_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_1209_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_1222_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_1234_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1247_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1259_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1272_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1284_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_2052_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1297_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1309_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1322_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1334_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1347_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1359_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1372_inst_req_0;
      RPIPE_maxpool_input_pipe_1555_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_1506_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_1967_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_2016_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_1998_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_2070_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_1519_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_1573_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_1627_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_1537_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_1591_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_2088_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_1980_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_1753_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_1609_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_2218_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_2034_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_1184_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_1197_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_1209_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_1222_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_1234_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_1247_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1259_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1272_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1284_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_2052_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1297_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1309_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1322_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1334_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1347_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1359_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1372_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_1555_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_1506_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_1967_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_2016_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_1998_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_2070_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_1519_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_1573_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_1627_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_1537_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_1591_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_2088_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_1980_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_1753_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_1609_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_2218_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_2034_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_1184_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_1197_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_1209_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_1222_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_1234_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1247_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1259_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1272_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1284_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_2052_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1297_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1309_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1322_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1334_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1347_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1359_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1372_inst_req_1;
      RPIPE_maxpool_input_pipe_1555_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_1506_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_1967_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_2016_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_1998_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_2070_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_1519_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_1573_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_1627_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_1537_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_1591_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_2088_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_1980_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_1753_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_1609_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_2218_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_2034_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_1184_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_1197_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_1209_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_1222_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_1234_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_1247_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1259_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1272_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1284_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_2052_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1297_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1309_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1322_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1334_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1347_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1359_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1372_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call105_1556 <= data_out(271 downto 264);
      call89_1507 <= data_out(263 downto 256);
      call164_1968 <= data_out(255 downto 248);
      call180_2017 <= data_out(247 downto 240);
      call174_1999 <= data_out(239 downto 232);
      call198_2071 <= data_out(231 downto 224);
      call93_1520 <= data_out(223 downto 216);
      call111_1574 <= data_out(215 downto 208);
      call129_1628 <= data_out(207 downto 200);
      call99_1538 <= data_out(199 downto 192);
      call117_1592 <= data_out(191 downto 184);
      call204_2089 <= data_out(183 downto 176);
      call168_1981 <= data_out(175 downto 168);
      callx_xi_1754 <= data_out(167 downto 160);
      call123_1610 <= data_out(159 downto 152);
      callx_xi359_2219 <= data_out(151 downto 144);
      call186_2035 <= data_out(143 downto 136);
      call_1185 <= data_out(135 downto 128);
      call2_1198 <= data_out(127 downto 120);
      call6_1210 <= data_out(119 downto 112);
      call11_1223 <= data_out(111 downto 104);
      call16_1235 <= data_out(103 downto 96);
      call21_1248 <= data_out(95 downto 88);
      call26_1260 <= data_out(87 downto 80);
      call31_1273 <= data_out(79 downto 72);
      call36_1285 <= data_out(71 downto 64);
      call192_2053 <= data_out(63 downto 56);
      call41_1298 <= data_out(55 downto 48);
      call46_1310 <= data_out(47 downto 40);
      call51_1323 <= data_out(39 downto 32);
      call56_1335 <= data_out(31 downto 24);
      call61_1348 <= data_out(23 downto 16);
      call66_1360 <= data_out(15 downto 8);
      call71_1373 <= data_out(7 downto 0);
      maxpool_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_1_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_1", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_2535_inst WPIPE_maxpool_output_pipe_2538_inst WPIPE_maxpool_output_pipe_2541_inst WPIPE_maxpool_output_pipe_2544_inst WPIPE_maxpool_output_pipe_2547_inst WPIPE_maxpool_output_pipe_2550_inst WPIPE_maxpool_output_pipe_2553_inst WPIPE_maxpool_output_pipe_2556_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_2535_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_2538_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_2541_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_2544_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_2547_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_2550_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2553_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2556_inst_req_0;
      WPIPE_maxpool_output_pipe_2535_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_2538_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_2541_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_2544_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_2547_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_2550_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_2553_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2556_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_2535_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_2538_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_2541_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_2544_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_2547_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_2550_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2553_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2556_inst_req_1;
      WPIPE_maxpool_output_pipe_2535_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_2538_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_2541_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_2544_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_2547_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_2550_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_2553_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2556_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv334_2534 & conv328_2524 & conv322_2514 & conv316_2504 & conv310_2494 & conv304_2484 & conv298_2474 & conv292_2464;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_num_out_pipe_2363_inst WPIPE_num_out_pipe_2366_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_num_out_pipe_2363_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_2366_inst_req_0;
      WPIPE_num_out_pipe_2363_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_num_out_pipe_2366_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_num_out_pipe_2363_inst_req_1;
      update_req_unguarded(0) <= WPIPE_num_out_pipe_2366_inst_req_1;
      WPIPE_num_out_pipe_2363_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_num_out_pipe_2366_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= add33_1282 & add43_1307;
      num_out_pipe_write_1_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_output_pipe_2308_inst WPIPE_output_pipe_2311_inst WPIPE_output_pipe_2314_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal sample_req, sample_ack : BooleanArray( 2 downto 0);
      signal update_req, update_ack : BooleanArray( 2 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 2 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      sample_req_unguarded(2) <= WPIPE_output_pipe_2308_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_output_pipe_2311_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_output_pipe_2314_inst_req_0;
      WPIPE_output_pipe_2308_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_output_pipe_2311_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_output_pipe_2314_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(2) <= WPIPE_output_pipe_2308_inst_req_1;
      update_req_unguarded(1) <= WPIPE_output_pipe_2311_inst_req_1;
      update_req_unguarded(0) <= WPIPE_output_pipe_2314_inst_req_1;
      WPIPE_output_pipe_2308_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_output_pipe_2311_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_output_pipe_2314_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      data_in <= add33_1282 & add43_1307 & add53_1332;
      output_pipe_write_2_gI: SplitGuardInterface generic map(name => "output_pipe_write_2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 3, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_2307_call call_stmt_2414_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_2307_call_req_0;
      reqL_unguarded(0) <= call_stmt_2414_call_req_0;
      call_stmt_2307_call_ack_0 <= ackL_unguarded(1);
      call_stmt_2414_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_2307_call_req_1;
      reqR_unguarded(0) <= call_stmt_2414_call_req_1;
      call_stmt_2307_call_ack_1 <= ackR_unguarded(1);
      call_stmt_2414_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call229_2307 <= data_out(127 downto 64);
      call275_2414 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2377_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2377_call_req_0;
      call_stmt_2377_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2377_call_req_1;
      call_stmt_2377_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv254_2374 & add23_1257;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(79 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2381_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2381_call_req_0;
      call_stmt_2381_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2381_call_req_1;
      call_stmt_2381_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add33_1282 & add23_1257 & add13_1232;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 48,
        owidth => 48,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(47 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_2459_call 
    sendB_call_group_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2459_call_req_0;
      call_stmt_2459_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2459_call_req_1;
      call_stmt_2459_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_3_gI: SplitGuardInterface generic map(name => "sendB_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv288_2457;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(63 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe4_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe4_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_6526_start: Boolean;
  signal convolve_CP_6526_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nacc1_2995_2595_buf_req_0 : boolean;
  signal phi_stmt_2596_req_0 : boolean;
  signal SUB_u16_u16_2586_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_2584_inst_ack_0 : boolean;
  signal nacc2_3004_2600_buf_ack_1 : boolean;
  signal phi_stmt_2596_req_1 : boolean;
  signal n_row_2986_2605_buf_req_1 : boolean;
  signal n_row_2986_2605_buf_ack_0 : boolean;
  signal phi_stmt_2601_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2784_inst_req_1 : boolean;
  signal W_store_kernel_2833_delayed_1_0_2935_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_2768_inst_req_1 : boolean;
  signal nacc1_2995_2595_buf_ack_1 : boolean;
  signal SUB_u16_u16_2581_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2734_inst_req_0 : boolean;
  signal phi_stmt_2590_ack_0 : boolean;
  signal SUB_u16_u16_2581_inst_req_1 : boolean;
  signal SUB_u16_u16_2586_inst_req_0 : boolean;
  signal n_row_2986_2605_buf_req_0 : boolean;
  signal phi_stmt_2606_req_1 : boolean;
  signal RPIPE_size_pipe_2584_inst_ack_1 : boolean;
  signal W_write_input_2652_delayed_1_0_2730_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe2_2768_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2784_inst_ack_1 : boolean;
  signal W_acc2_2781_delayed_1_0_2873_inst_req_0 : boolean;
  signal W_write_input_2652_delayed_1_0_2730_inst_req_1 : boolean;
  signal W_acc2_2781_delayed_1_0_2873_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_2584_inst_req_0 : boolean;
  signal nacc2_3004_2600_buf_req_0 : boolean;
  signal nacc2_3004_2600_buf_ack_0 : boolean;
  signal phi_stmt_2606_ack_0 : boolean;
  signal phi_stmt_2590_req_1 : boolean;
  signal W_read_k_2718_delayed_1_0_2804_inst_ack_1 : boolean;
  signal n_row_2986_2605_buf_ack_1 : boolean;
  signal SUB_u16_u16_2586_inst_req_1 : boolean;
  signal W_write_input_2652_delayed_1_0_2730_inst_ack_0 : boolean;
  signal n_col_2978_2610_buf_ack_0 : boolean;
  signal do_while_stmt_2588_branch_req_0 : boolean;
  signal SUB_u16_u16_2586_inst_ack_1 : boolean;
  signal W_store_kernel_2833_delayed_1_0_2935_inst_req_0 : boolean;
  signal n_col_2978_2610_buf_req_1 : boolean;
  signal W_read_k_2718_delayed_1_0_2804_inst_req_1 : boolean;
  signal n_col_2978_2610_buf_ack_1 : boolean;
  signal phi_stmt_2601_ack_0 : boolean;
  signal phi_stmt_2590_req_0 : boolean;
  signal nacc1_2995_2595_buf_ack_0 : boolean;
  signal n_col_2978_2610_buf_req_0 : boolean;
  signal phi_stmt_2606_req_0 : boolean;
  signal phi_stmt_2596_ack_0 : boolean;
  signal nacc1_2995_2595_buf_req_1 : boolean;
  signal nacc2_3004_2600_buf_req_1 : boolean;
  signal phi_stmt_2601_req_1 : boolean;
  signal RPIPE_size_pipe_2584_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2734_inst_ack_0 : boolean;
  signal W_num_done_2880_delayed_1_0_2987_inst_ack_1 : boolean;
  signal W_num_done_2886_delayed_1_0_2996_inst_req_0 : boolean;
  signal W_num_done_2886_delayed_1_0_2996_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe3_2772_inst_req_0 : boolean;
  signal W_acc2_2781_delayed_1_0_2873_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe3_2772_inst_ack_0 : boolean;
  signal W_acc2_2781_delayed_1_0_2873_inst_ack_1 : boolean;
  signal W_store_kernel_2837_delayed_1_0_2942_inst_req_1 : boolean;
  signal W_write_input_2648_delayed_1_0_2723_inst_req_0 : boolean;
  signal W_store_kernel_2833_delayed_1_0_2935_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe3_2772_inst_req_1 : boolean;
  signal W_store_kernel_2829_delayed_1_0_2928_inst_req_0 : boolean;
  signal W_store_kernel_2833_delayed_1_0_2935_inst_ack_1 : boolean;
  signal RPIPE_num_out_pipe_2574_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_2574_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2574_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_2574_inst_ack_1 : boolean;
  signal SUB_u16_u16_2576_inst_req_0 : boolean;
  signal SUB_u16_u16_2576_inst_ack_0 : boolean;
  signal SUB_u16_u16_2576_inst_req_1 : boolean;
  signal SUB_u16_u16_2576_inst_ack_1 : boolean;
  signal RPIPE_num_out_pipe_2579_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_2579_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_2579_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_2579_inst_ack_1 : boolean;
  signal SUB_u16_u16_2581_inst_req_0 : boolean;
  signal SUB_u16_u16_2581_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2727_inst_ack_1 : boolean;
  signal phi_stmt_2611_req_1 : boolean;
  signal phi_stmt_2611_req_0 : boolean;
  signal phi_stmt_2611_ack_0 : boolean;
  signal n_num_2967_2616_buf_req_0 : boolean;
  signal n_num_2967_2616_buf_ack_0 : boolean;
  signal n_num_2967_2616_buf_req_1 : boolean;
  signal n_num_2967_2616_buf_ack_1 : boolean;
  signal phi_stmt_2617_req_1 : boolean;
  signal phi_stmt_2617_req_0 : boolean;
  signal phi_stmt_2617_ack_0 : boolean;
  signal W_read_k_2718_delayed_1_0_2804_inst_ack_0 : boolean;
  signal W_num_done_2880_delayed_1_0_2987_inst_req_1 : boolean;
  signal W_store_kernel_2837_delayed_1_0_2942_inst_ack_0 : boolean;
  signal W_read_k_2718_delayed_1_0_2804_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe2_2768_inst_ack_0 : boolean;
  signal n_chl_2956_2621_buf_req_0 : boolean;
  signal n_chl_2956_2621_buf_ack_0 : boolean;
  signal W_write_input_2652_delayed_1_0_2730_inst_req_0 : boolean;
  signal n_chl_2956_2621_buf_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2784_inst_ack_0 : boolean;
  signal n_chl_2956_2621_buf_ack_1 : boolean;
  signal RPIPE_kernel_pipe2_2768_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_2634_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2784_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_2634_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_2634_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_2634_inst_ack_1 : boolean;
  signal W_store_kernel_2837_delayed_1_0_2942_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2720_inst_ack_1 : boolean;
  signal RPIPE_input_pipe2_2638_inst_req_0 : boolean;
  signal RPIPE_input_pipe2_2638_inst_ack_0 : boolean;
  signal RPIPE_input_pipe2_2638_inst_req_1 : boolean;
  signal RPIPE_input_pipe2_2638_inst_ack_1 : boolean;
  signal SUB_u16_u16_2910_inst_ack_1 : boolean;
  signal W_read_k_2712_delayed_1_0_2795_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_2764_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2720_inst_req_1 : boolean;
  signal RPIPE_input_pipe3_2642_inst_req_0 : boolean;
  signal RPIPE_input_pipe3_2642_inst_ack_0 : boolean;
  signal RPIPE_input_pipe3_2642_inst_req_1 : boolean;
  signal RPIPE_input_pipe3_2642_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2939_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2939_inst_req_1 : boolean;
  signal SUB_u16_u16_2910_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_2764_inst_req_1 : boolean;
  signal W_read_k_2712_delayed_1_0_2795_inst_req_1 : boolean;
  signal RPIPE_input_pipe4_2646_inst_req_0 : boolean;
  signal RPIPE_input_pipe4_2646_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2780_inst_ack_1 : boolean;
  signal RPIPE_input_pipe4_2646_inst_req_1 : boolean;
  signal RPIPE_input_pipe4_2646_inst_ack_1 : boolean;
  signal W_write_input_2648_delayed_1_0_2723_inst_ack_1 : boolean;
  signal W_write_input_2648_delayed_1_0_2723_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2780_inst_req_1 : boolean;
  signal W_write_input_2648_delayed_1_0_2723_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2650_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2650_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2650_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_2650_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2939_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_2764_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_2764_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2946_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2654_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2780_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2654_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2654_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2780_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_2654_inst_ack_1 : boolean;
  signal SUB_u16_u16_2910_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2939_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2932_inst_ack_1 : boolean;
  signal SUB_u16_u16_2910_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2946_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2658_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2658_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2727_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2658_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_2658_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2932_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2662_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2662_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2662_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_2662_inst_ack_1 : boolean;
  signal W_read_k_2712_delayed_1_0_2795_inst_ack_0 : boolean;
  signal W_read_k_2712_delayed_1_0_2795_inst_req_0 : boolean;
  signal W_read_ip_2608_delayed_1_0_2664_inst_req_0 : boolean;
  signal W_read_ip_2608_delayed_1_0_2664_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2932_inst_ack_0 : boolean;
  signal W_read_ip_2608_delayed_1_0_2664_inst_req_1 : boolean;
  signal W_read_ip_2608_delayed_1_0_2664_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2932_inst_req_0 : boolean;
  signal W_read_ip_2614_delayed_1_0_2673_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2776_inst_ack_1 : boolean;
  signal W_read_ip_2614_delayed_1_0_2673_inst_ack_0 : boolean;
  signal W_read_ip_2614_delayed_1_0_2673_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2776_inst_req_1 : boolean;
  signal W_read_ip_2614_delayed_1_0_2673_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2946_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2734_inst_ack_1 : boolean;
  signal W_read_ip_2620_delayed_1_0_2682_inst_req_0 : boolean;
  signal W_read_ip_2620_delayed_1_0_2682_inst_ack_0 : boolean;
  signal W_read_ip_2620_delayed_1_0_2682_inst_req_1 : boolean;
  signal W_read_ip_2620_delayed_1_0_2682_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2734_inst_req_1 : boolean;
  signal W_read_ip_2626_delayed_1_0_2691_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2776_inst_ack_0 : boolean;
  signal W_read_ip_2626_delayed_1_0_2691_inst_ack_0 : boolean;
  signal W_read_ip_2626_delayed_1_0_2691_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2776_inst_req_0 : boolean;
  signal W_read_ip_2626_delayed_1_0_2691_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2946_inst_req_0 : boolean;
  signal W_read_k_2706_delayed_1_0_2786_inst_ack_1 : boolean;
  signal W_read_k_2706_delayed_1_0_2786_inst_req_1 : boolean;
  signal W_write_input_2640_delayed_1_0_2709_inst_req_0 : boolean;
  signal W_write_input_2640_delayed_1_0_2709_inst_ack_0 : boolean;
  signal W_store_kernel_2829_delayed_1_0_2928_inst_ack_1 : boolean;
  signal W_write_input_2640_delayed_1_0_2709_inst_req_1 : boolean;
  signal W_write_input_2640_delayed_1_0_2709_inst_ack_1 : boolean;
  signal W_acc1_2772_delayed_1_0_2861_inst_ack_1 : boolean;
  signal W_acc1_2772_delayed_1_0_2861_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2727_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2713_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2713_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2727_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2713_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2713_inst_ack_1 : boolean;
  signal W_store_kernel_2829_delayed_1_0_2928_inst_req_1 : boolean;
  signal W_num_done_2880_delayed_1_0_2987_inst_ack_0 : boolean;
  signal W_read_k_2706_delayed_1_0_2786_inst_ack_0 : boolean;
  signal W_write_input_2644_delayed_1_0_2716_inst_req_0 : boolean;
  signal W_write_input_2644_delayed_1_0_2716_inst_ack_0 : boolean;
  signal W_store_kernel_2829_delayed_1_0_2928_inst_ack_0 : boolean;
  signal W_write_input_2644_delayed_1_0_2716_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe3_2772_inst_ack_1 : boolean;
  signal W_write_input_2644_delayed_1_0_2716_inst_ack_1 : boolean;
  signal W_store_kernel_2837_delayed_1_0_2942_inst_ack_1 : boolean;
  signal W_read_k_2706_delayed_1_0_2786_inst_req_0 : boolean;
  signal W_num_done_2880_delayed_1_0_2987_inst_req_0 : boolean;
  signal W_acc1_2772_delayed_1_0_2861_inst_ack_0 : boolean;
  signal W_acc1_2772_delayed_1_0_2861_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2720_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2720_inst_ack_0 : boolean;
  signal W_num_done_2886_delayed_1_0_2996_inst_req_1 : boolean;
  signal W_num_done_2886_delayed_1_0_2996_inst_ack_1 : boolean;
  signal W_num_done_2891_delayed_1_0_3005_inst_req_0 : boolean;
  signal W_num_done_2891_delayed_1_0_3005_inst_ack_0 : boolean;
  signal W_num_done_2891_delayed_1_0_3005_inst_req_1 : boolean;
  signal W_num_done_2891_delayed_1_0_3005_inst_ack_1 : boolean;
  signal type_cast_3011_inst_req_0 : boolean;
  signal type_cast_3011_inst_ack_0 : boolean;
  signal type_cast_3011_inst_req_1 : boolean;
  signal type_cast_3011_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_3009_inst_req_0 : boolean;
  signal WPIPE_output_pipe_3009_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_3009_inst_req_1 : boolean;
  signal WPIPE_output_pipe_3009_inst_ack_1 : boolean;
  signal W_num_done_2896_delayed_1_0_3013_inst_req_0 : boolean;
  signal W_num_done_2896_delayed_1_0_3013_inst_ack_0 : boolean;
  signal W_num_done_2896_delayed_1_0_3013_inst_req_1 : boolean;
  signal W_num_done_2896_delayed_1_0_3013_inst_ack_1 : boolean;
  signal type_cast_3019_inst_req_0 : boolean;
  signal type_cast_3019_inst_ack_0 : boolean;
  signal type_cast_3019_inst_req_1 : boolean;
  signal type_cast_3019_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_3017_inst_req_0 : boolean;
  signal WPIPE_output_pipe_3017_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_3017_inst_req_1 : boolean;
  signal WPIPE_output_pipe_3017_inst_ack_1 : boolean;
  signal do_while_stmt_2588_branch_ack_0 : boolean;
  signal do_while_stmt_2588_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3024_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3024_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_3024_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_3024_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_6526_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_6526_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_6526_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_6526_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_6526: Block -- control-path 
    signal convolve_CP_6526_elements: BooleanArray(323 downto 0);
    -- 
  begin -- 
    convolve_CP_6526_elements(0) <= convolve_CP_6526_start;
    convolve_CP_6526_symbol <= convolve_CP_6526_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	323 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2571/$entry
      -- CP-element group 0: 	 branch_block_stmt_2571/branch_block_stmt_2571__entry__
      -- CP-element group 0: 	 branch_block_stmt_2571/merge_stmt_2572__entry__
      -- CP-element group 0: 	 branch_block_stmt_2571/merge_stmt_2572_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_2571/merge_stmt_2572__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_2571/merge_stmt_2572__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2571/$exit
      -- CP-element group 1: 	 branch_block_stmt_2571/branch_block_stmt_2571__exit__
      -- 
    convolve_CP_6526_elements(1) <= false; 
    -- CP-element group 2:  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	320 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	321 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2571/do_while_stmt_2588__exit__
      -- CP-element group 2: 	 branch_block_stmt_2571/assign_stmt_3026__entry__
      -- CP-element group 2: 	 branch_block_stmt_2571/assign_stmt_3026/$entry
      -- CP-element group 2: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_Sample/req
      -- 
    req_7578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(2), ack => WPIPE_input_done_pipe_3024_inst_req_0); -- 
    convolve_CP_6526_elements(2) <= convolve_CP_6526_elements(320);
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	323 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_update_start_
      -- CP-element group 3: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_Update/cr
      -- 
    ra_6558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2574_inst_ack_0, ack => convolve_CP_6526_elements(3)); -- 
    cr_6562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(3), ack => RPIPE_num_out_pipe_2574_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_Sample/rr
      -- 
    ca_6563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2574_inst_ack_1, ack => convolve_CP_6526_elements(4)); -- 
    rr_6567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(4), ack => SUB_u16_u16_2576_inst_req_0); -- 
    rr_6585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(4), ack => RPIPE_num_out_pipe_2579_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_Sample/ra
      -- 
    ra_6568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2576_inst_ack_0, ack => convolve_CP_6526_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	323 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	15 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_Update/ca
      -- 
    ca_6573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2576_inst_ack_1, ack => convolve_CP_6526_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_update_start_
      -- CP-element group 7: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_Update/cr
      -- 
    ra_6586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2579_inst_ack_0, ack => convolve_CP_6526_elements(7)); -- 
    cr_6590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(7), ack => RPIPE_num_out_pipe_2579_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2579_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_Sample/rr
      -- 
    ca_6591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_2579_inst_ack_1, ack => convolve_CP_6526_elements(8)); -- 
    rr_6595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(8), ack => SUB_u16_u16_2581_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_Sample/ra
      -- 
    ra_6596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2581_inst_ack_0, ack => convolve_CP_6526_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	323 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_update_completed_
      -- 
    ca_6601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2581_inst_ack_1, ack => convolve_CP_6526_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	323 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_update_start_
      -- CP-element group 11: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_Update/cr
      -- 
    ra_6614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_2584_inst_ack_0, ack => convolve_CP_6526_elements(11)); -- 
    cr_6618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(11), ack => RPIPE_size_pipe_2584_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_Update/$exit
      -- 
    ca_6619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_2584_inst_ack_1, ack => convolve_CP_6526_elements(12)); -- 
    rr_6623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(12), ack => SUB_u16_u16_2586_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_Sample/$exit
      -- 
    ra_6624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2586_inst_ack_0, ack => convolve_CP_6526_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	323 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_Update/ca
      -- 
    ca_6629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2586_inst_ack_1, ack => convolve_CP_6526_elements(14)); -- 
    -- CP-element group 15:  join  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	6 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587__exit__
      -- CP-element group 15: 	 branch_block_stmt_2571/do_while_stmt_2588__entry__
      -- CP-element group 15: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/$exit
      -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(6) & convolve_CP_6526_elements(10) & convolve_CP_6526_elements(14);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588__entry__
      -- CP-element group 16: 	 branch_block_stmt_2571/do_while_stmt_2588/$entry
      -- 
    convolve_CP_6526_elements(16) <= convolve_CP_6526_elements(15);
    -- CP-element group 17:  merge  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	320 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588__exit__
      -- 
    -- Element group convolve_CP_6526_elements(17) is bound as output of CP function.
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2571/do_while_stmt_2588/loop_back
      -- 
    -- Element group convolve_CP_6526_elements(18) is bound as output of CP function.
    -- CP-element group 19:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	318 
    -- CP-element group 19: 	319 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2571/do_while_stmt_2588/condition_done
      -- CP-element group 19: 	 branch_block_stmt_2571/do_while_stmt_2588/loop_exit/$entry
      -- CP-element group 19: 	 branch_block_stmt_2571/do_while_stmt_2588/loop_taken/$entry
      -- 
    convolve_CP_6526_elements(19) <= convolve_CP_6526_elements(24);
    -- CP-element group 20:  branch  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	317 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2571/do_while_stmt_2588/loop_body_done
      -- 
    convolve_CP_6526_elements(20) <= convolve_CP_6526_elements(317);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	109 
    -- CP-element group 21: 	35 
    -- CP-element group 21: 	54 
    -- CP-element group 21: 	73 
    -- CP-element group 21: 	92 
    -- CP-element group 21: 	128 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_6526_elements(21) <= convolve_CP_6526_elements(18);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	111 
    -- CP-element group 22: 	37 
    -- CP-element group 22: 	56 
    -- CP-element group 22: 	75 
    -- CP-element group 22: 	94 
    -- CP-element group 22: 	130 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_6526_elements(22) <= convolve_CP_6526_elements(16);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	225 
    -- CP-element group 23: 	217 
    -- CP-element group 23: 	221 
    -- CP-element group 23: 	105 
    -- CP-element group 23: 	106 
    -- CP-element group 23: 	237 
    -- CP-element group 23: 	229 
    -- CP-element group 23: 	233 
    -- CP-element group 23: 	261 
    -- CP-element group 23: 	29 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	48 
    -- CP-element group 23: 	49 
    -- CP-element group 23: 	316 
    -- CP-element group 23: 	67 
    -- CP-element group 23: 	68 
    -- CP-element group 23: 	86 
    -- CP-element group 23: 	87 
    -- CP-element group 23: 	169 
    -- CP-element group 23: 	122 
    -- CP-element group 23: 	123 
    -- CP-element group 23: 	149 
    -- CP-element group 23: 	153 
    -- CP-element group 23: 	157 
    -- CP-element group 23: 	161 
    -- CP-element group 23: 	165 
    -- CP-element group 23: 	141 
    -- CP-element group 23: 	145 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/$entry
      -- CP-element group 23: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_6526_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	108 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	316 
    -- CP-element group 24: 	72 
    -- CP-element group 24: 	91 
    -- CP-element group 24: 	127 
    -- CP-element group 24: 	264 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/condition_evaluated
      -- 
    condition_evaluated_6644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(24), ack => do_while_stmt_2588_branch_req_0); -- 
    convolve_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(28) & convolve_CP_6526_elements(316) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(127) & convolve_CP_6526_elements(264);
      gj_convolve_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	105 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	48 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	86 
    -- CP-element group 25: 	122 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	31 
    -- CP-element group 25: 	50 
    -- CP-element group 25: 	69 
    -- CP-element group 25: 	88 
    -- CP-element group 25: 	124 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/aggregated_phi_sample_req
      -- CP-element group 25: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_sample_start__ps
      -- 
    convolve_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(105) & convolve_CP_6526_elements(29) & convolve_CP_6526_elements(48) & convolve_CP_6526_elements(67) & convolve_CP_6526_elements(86) & convolve_CP_6526_elements(122) & convolve_CP_6526_elements(28);
      gj_convolve_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	107 
    -- CP-element group 26: 	32 
    -- CP-element group 26: 	51 
    -- CP-element group 26: 	70 
    -- CP-element group 26: 	89 
    -- CP-element group 26: 	125 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	287 
    -- CP-element group 26: 	222 
    -- CP-element group 26: 	226 
    -- CP-element group 26: 	218 
    -- CP-element group 26: 	242 
    -- CP-element group 26: 	246 
    -- CP-element group 26: 	250 
    -- CP-element group 26: 	254 
    -- CP-element group 26: 	238 
    -- CP-element group 26: 	230 
    -- CP-element group 26: 	234 
    -- CP-element group 26: 	258 
    -- CP-element group 26: 	291 
    -- CP-element group 26: 	317 
    -- CP-element group 26: 	174 
    -- CP-element group 26: 	178 
    -- CP-element group 26: 	166 
    -- CP-element group 26: 	170 
    -- CP-element group 26: 	146 
    -- CP-element group 26: 	150 
    -- CP-element group 26: 	154 
    -- CP-element group 26: 	158 
    -- CP-element group 26: 	162 
    -- CP-element group 26: 	142 
    -- CP-element group 26: 	182 
    -- CP-element group 26: 	186 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	105 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	48 
    -- CP-element group 26: 	67 
    -- CP-element group 26: 	86 
    -- CP-element group 26: 	122 
    -- CP-element group 26:  members (7) 
      -- CP-element group 26: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/aggregated_phi_sample_ack
      -- CP-element group 26: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_sample_completed_
      -- 
    convolve_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(107) & convolve_CP_6526_elements(32) & convolve_CP_6526_elements(51) & convolve_CP_6526_elements(70) & convolve_CP_6526_elements(89) & convolve_CP_6526_elements(125);
      gj_convolve_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	106 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	49 
    -- CP-element group 27: 	68 
    -- CP-element group 27: 	87 
    -- CP-element group 27: 	123 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	33 
    -- CP-element group 27: 	52 
    -- CP-element group 27: 	71 
    -- CP-element group 27: 	90 
    -- CP-element group 27: 	126 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/aggregated_phi_update_req
      -- CP-element group 27: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_update_start__ps
      -- 
    convolve_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(106) & convolve_CP_6526_elements(30) & convolve_CP_6526_elements(49) & convolve_CP_6526_elements(68) & convolve_CP_6526_elements(87) & convolve_CP_6526_elements(123);
      gj_convolve_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	108 
    -- CP-element group 28: 	34 
    -- CP-element group 28: 	53 
    -- CP-element group 28: 	72 
    -- CP-element group 28: 	91 
    -- CP-element group 28: 	127 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(34) & convolve_CP_6526_elements(53) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(127);
      gj_convolve_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	224 
    -- CP-element group 29: 	220 
    -- CP-element group 29: 	244 
    -- CP-element group 29: 	248 
    -- CP-element group 29: 	252 
    -- CP-element group 29: 	236 
    -- CP-element group 29: 	240 
    -- CP-element group 29: 	228 
    -- CP-element group 29: 	232 
    -- CP-element group 29: 	256 
    -- CP-element group 29: 	289 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	176 
    -- CP-element group 29: 	168 
    -- CP-element group 29: 	148 
    -- CP-element group 29: 	152 
    -- CP-element group 29: 	160 
    -- CP-element group 29: 	164 
    -- CP-element group 29: 	144 
    -- CP-element group 29: 	180 
    -- CP-element group 29: 	184 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_sample_start_
      -- 
    convolve_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(224) & convolve_CP_6526_elements(220) & convolve_CP_6526_elements(244) & convolve_CP_6526_elements(248) & convolve_CP_6526_elements(252) & convolve_CP_6526_elements(236) & convolve_CP_6526_elements(240) & convolve_CP_6526_elements(228) & convolve_CP_6526_elements(232) & convolve_CP_6526_elements(256) & convolve_CP_6526_elements(289) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(176) & convolve_CP_6526_elements(168) & convolve_CP_6526_elements(148) & convolve_CP_6526_elements(152) & convolve_CP_6526_elements(160) & convolve_CP_6526_elements(164) & convolve_CP_6526_elements(144) & convolve_CP_6526_elements(180) & convolve_CP_6526_elements(184);
      gj_convolve_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	255 
    -- CP-element group 30: 	34 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	27 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_update_start_
      -- 
    convolve_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(255) & convolve_CP_6526_elements(34);
      gj_convolve_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	25 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_sample_start__ps
      -- 
    convolve_CP_6526_elements(31) <= convolve_CP_6526_elements(25);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	26 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_sample_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(32) is bound as output of CP function.
    -- CP-element group 33:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	27 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_update_start__ps
      -- 
    convolve_CP_6526_elements(33) <= convolve_CP_6526_elements(27);
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	253 
    -- CP-element group 34: 	28 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	30 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_update_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(34) is bound as output of CP function.
    -- CP-element group 35:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	21 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_loopback_trigger
      -- 
    convolve_CP_6526_elements(35) <= convolve_CP_6526_elements(21);
    -- CP-element group 36:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_loopback_sample_req
      -- CP-element group 36: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_loopback_sample_req_ps
      -- 
    phi_stmt_2590_loopback_sample_req_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2590_loopback_sample_req_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(36), ack => phi_stmt_2590_req_1); -- 
    -- Element group convolve_CP_6526_elements(36) is bound as output of CP function.
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	22 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_entry_trigger
      -- 
    convolve_CP_6526_elements(37) <= convolve_CP_6526_elements(22);
    -- CP-element group 38:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_entry_sample_req_ps
      -- CP-element group 38: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_entry_sample_req
      -- 
    phi_stmt_2590_entry_sample_req_6662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2590_entry_sample_req_6662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(38), ack => phi_stmt_2590_req_0); -- 
    -- Element group convolve_CP_6526_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_phi_mux_ack_ps
      -- CP-element group 39: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2590_phi_mux_ack
      -- 
    phi_stmt_2590_phi_mux_ack_6665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2590_ack_0, ack => convolve_CP_6526_elements(39)); -- 
    -- CP-element group 40:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2594_sample_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2594_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2594_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2594_sample_start__ps
      -- 
    -- Element group convolve_CP_6526_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2594_update_start__ps
      -- CP-element group 41: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2594_update_start_
      -- 
    -- Element group convolve_CP_6526_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2594_update_completed__ps
      -- 
    convolve_CP_6526_elements(42) <= convolve_CP_6526_elements(43);
    -- CP-element group 43:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	42 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2594_update_completed_
      -- 
    -- Element group convolve_CP_6526_elements(43) is a control-delay.
    cp_element_43_delay: control_delay_element  generic map(name => " 43_delay", delay_value => 1)  port map(req => convolve_CP_6526_elements(41), ack => convolve_CP_6526_elements(43), clk => clk, reset =>reset);
    -- CP-element group 44:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_Sample/req
      -- CP-element group 44: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_sample_start__ps
      -- CP-element group 44: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_sample_start_
      -- 
    req_6686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(44), ack => nacc1_2995_2595_buf_req_0); -- 
    -- Element group convolve_CP_6526_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_update_start__ps
      -- CP-element group 45: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_Update/req
      -- CP-element group 45: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_update_start_
      -- 
    req_6691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(45), ack => nacc1_2995_2595_buf_req_1); -- 
    -- Element group convolve_CP_6526_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_sample_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_sample_completed_
      -- 
    ack_6687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc1_2995_2595_buf_ack_0, ack => convolve_CP_6526_elements(46)); -- 
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_update_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc1_2595_Update/$exit
      -- 
    ack_6692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc1_2995_2595_buf_ack_1, ack => convolve_CP_6526_elements(47)); -- 
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	23 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	224 
    -- CP-element group 48: 	220 
    -- CP-element group 48: 	244 
    -- CP-element group 48: 	248 
    -- CP-element group 48: 	252 
    -- CP-element group 48: 	236 
    -- CP-element group 48: 	240 
    -- CP-element group 48: 	228 
    -- CP-element group 48: 	232 
    -- CP-element group 48: 	260 
    -- CP-element group 48: 	293 
    -- CP-element group 48: 	26 
    -- CP-element group 48: 	172 
    -- CP-element group 48: 	168 
    -- CP-element group 48: 	148 
    -- CP-element group 48: 	152 
    -- CP-element group 48: 	156 
    -- CP-element group 48: 	164 
    -- CP-element group 48: 	180 
    -- CP-element group 48: 	184 
    -- CP-element group 48: 	188 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	25 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_sample_start_
      -- 
    convolve_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(224) & convolve_CP_6526_elements(220) & convolve_CP_6526_elements(244) & convolve_CP_6526_elements(248) & convolve_CP_6526_elements(252) & convolve_CP_6526_elements(236) & convolve_CP_6526_elements(240) & convolve_CP_6526_elements(228) & convolve_CP_6526_elements(232) & convolve_CP_6526_elements(260) & convolve_CP_6526_elements(293) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(172) & convolve_CP_6526_elements(168) & convolve_CP_6526_elements(148) & convolve_CP_6526_elements(152) & convolve_CP_6526_elements(156) & convolve_CP_6526_elements(164) & convolve_CP_6526_elements(180) & convolve_CP_6526_elements(184) & convolve_CP_6526_elements(188);
      gj_convolve_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	23 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	259 
    -- CP-element group 49: 	53 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	27 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_update_start_
      -- 
    convolve_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(259) & convolve_CP_6526_elements(53);
      gj_convolve_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	25 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_sample_start__ps
      -- 
    convolve_CP_6526_elements(50) <= convolve_CP_6526_elements(25);
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	26 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_sample_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	27 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_update_start__ps
      -- 
    convolve_CP_6526_elements(52) <= convolve_CP_6526_elements(27);
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	257 
    -- CP-element group 53: 	28 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	49 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_update_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_update_completed_
      -- 
    -- Element group convolve_CP_6526_elements(53) is bound as output of CP function.
    -- CP-element group 54:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	21 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_loopback_trigger
      -- 
    convolve_CP_6526_elements(54) <= convolve_CP_6526_elements(21);
    -- CP-element group 55:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_loopback_sample_req
      -- CP-element group 55: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_loopback_sample_req_ps
      -- 
    phi_stmt_2596_loopback_sample_req_6703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2596_loopback_sample_req_6703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(55), ack => phi_stmt_2596_req_1); -- 
    -- Element group convolve_CP_6526_elements(55) is bound as output of CP function.
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	22 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_entry_trigger
      -- 
    convolve_CP_6526_elements(56) <= convolve_CP_6526_elements(22);
    -- CP-element group 57:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_entry_sample_req
      -- CP-element group 57: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_entry_sample_req_ps
      -- 
    phi_stmt_2596_entry_sample_req_6706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2596_entry_sample_req_6706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(57), ack => phi_stmt_2596_req_0); -- 
    -- Element group convolve_CP_6526_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_phi_mux_ack
      -- CP-element group 58: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2596_phi_mux_ack_ps
      -- 
    phi_stmt_2596_phi_mux_ack_6709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2596_ack_0, ack => convolve_CP_6526_elements(58)); -- 
    -- CP-element group 59:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2599_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2599_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2599_sample_start__ps
      -- CP-element group 59: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2599_sample_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(59) is bound as output of CP function.
    -- CP-element group 60:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2599_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2599_update_start__ps
      -- 
    -- Element group convolve_CP_6526_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2599_update_completed__ps
      -- 
    convolve_CP_6526_elements(61) <= convolve_CP_6526_elements(62);
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	61 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2599_update_completed_
      -- 
    -- Element group convolve_CP_6526_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => convolve_CP_6526_elements(60), ack => convolve_CP_6526_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_sample_start__ps
      -- CP-element group 63: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_sample_start_
      -- 
    req_6730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(63), ack => nacc2_3004_2600_buf_req_0); -- 
    -- Element group convolve_CP_6526_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_update_start_
      -- CP-element group 64: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_update_start__ps
      -- CP-element group 64: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_Update/req
      -- 
    req_6735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(64), ack => nacc2_3004_2600_buf_req_1); -- 
    -- Element group convolve_CP_6526_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_sample_completed__ps
      -- CP-element group 65: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_Sample/ack
      -- CP-element group 65: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_sample_completed_
      -- 
    ack_6731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc2_3004_2600_buf_ack_0, ack => convolve_CP_6526_elements(65)); -- 
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_Update/ack
      -- CP-element group 66: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_nacc2_2600_update_completed__ps
      -- 
    ack_6736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc2_3004_2600_buf_ack_1, ack => convolve_CP_6526_elements(66)); -- 
    -- CP-element group 67:  join  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	23 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	26 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	25 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_sample_start_
      -- 
    convolve_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(26);
      gj_convolve_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	23 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	281 
    -- CP-element group 68: 	222 
    -- CP-element group 68: 	226 
    -- CP-element group 68: 	274 
    -- CP-element group 68: 	218 
    -- CP-element group 68: 	243 
    -- CP-element group 68: 	247 
    -- CP-element group 68: 	251 
    -- CP-element group 68: 	238 
    -- CP-element group 68: 	230 
    -- CP-element group 68: 	234 
    -- CP-element group 68: 	72 
    -- CP-element group 68: 	267 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	27 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_update_start_
      -- 
    convolve_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(281) & convolve_CP_6526_elements(222) & convolve_CP_6526_elements(226) & convolve_CP_6526_elements(274) & convolve_CP_6526_elements(218) & convolve_CP_6526_elements(243) & convolve_CP_6526_elements(247) & convolve_CP_6526_elements(251) & convolve_CP_6526_elements(238) & convolve_CP_6526_elements(230) & convolve_CP_6526_elements(234) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(267);
      gj_convolve_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	25 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_sample_start__ps
      -- 
    convolve_CP_6526_elements(69) <= convolve_CP_6526_elements(25);
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	26 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_sample_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(70) is bound as output of CP function.
    -- CP-element group 71:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	27 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_update_start__ps
      -- 
    convolve_CP_6526_elements(71) <= convolve_CP_6526_elements(27);
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	222 
    -- CP-element group 72: 	226 
    -- CP-element group 72: 	272 
    -- CP-element group 72: 	279 
    -- CP-element group 72: 	218 
    -- CP-element group 72: 	245 
    -- CP-element group 72: 	249 
    -- CP-element group 72: 	238 
    -- CP-element group 72: 	241 
    -- CP-element group 72: 	230 
    -- CP-element group 72: 	234 
    -- CP-element group 72: 	24 
    -- CP-element group 72: 	28 
    -- CP-element group 72: 	265 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	68 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_update_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(72) is bound as output of CP function.
    -- CP-element group 73:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	21 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_loopback_trigger
      -- 
    convolve_CP_6526_elements(73) <= convolve_CP_6526_elements(21);
    -- CP-element group 74:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_loopback_sample_req_ps
      -- CP-element group 74: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_loopback_sample_req
      -- 
    phi_stmt_2601_loopback_sample_req_6747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2601_loopback_sample_req_6747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(74), ack => phi_stmt_2601_req_1); -- 
    -- Element group convolve_CP_6526_elements(74) is bound as output of CP function.
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	22 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_entry_trigger
      -- 
    convolve_CP_6526_elements(75) <= convolve_CP_6526_elements(22);
    -- CP-element group 76:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_entry_sample_req_ps
      -- CP-element group 76: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_entry_sample_req
      -- 
    phi_stmt_2601_entry_sample_req_6750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2601_entry_sample_req_6750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(76), ack => phi_stmt_2601_req_0); -- 
    -- Element group convolve_CP_6526_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_phi_mux_ack_ps
      -- CP-element group 77: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2601_phi_mux_ack
      -- 
    phi_stmt_2601_phi_mux_ack_6753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2601_ack_0, ack => convolve_CP_6526_elements(77)); -- 
    -- CP-element group 78:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (4) 
      -- CP-element group 78: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2604_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2604_sample_completed__ps
      -- CP-element group 78: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2604_sample_start__ps
      -- CP-element group 78: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2604_sample_start_
      -- 
    -- Element group convolve_CP_6526_elements(78) is bound as output of CP function.
    -- CP-element group 79:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2604_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2604_update_start__ps
      -- 
    -- Element group convolve_CP_6526_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2604_update_completed__ps
      -- 
    convolve_CP_6526_elements(80) <= convolve_CP_6526_elements(81);
    -- CP-element group 81:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	80 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2604_update_completed_
      -- 
    -- Element group convolve_CP_6526_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convolve_CP_6526_elements(79), ack => convolve_CP_6526_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_Sample/req
      -- CP-element group 82: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_sample_start__ps
      -- CP-element group 82: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_Sample/$entry
      -- 
    req_6774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(82), ack => n_row_2986_2605_buf_req_0); -- 
    -- Element group convolve_CP_6526_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_Update/req
      -- CP-element group 83: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_update_start__ps
      -- CP-element group 83: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_update_start_
      -- 
    req_6779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(83), ack => n_row_2986_2605_buf_req_1); -- 
    -- Element group convolve_CP_6526_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_Sample/ack
      -- CP-element group 84: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_sample_completed__ps
      -- CP-element group 84: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_Sample/$exit
      -- 
    ack_6775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_2986_2605_buf_ack_0, ack => convolve_CP_6526_elements(84)); -- 
    -- CP-element group 85:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_update_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_row_2605_update_completed_
      -- 
    ack_6780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_2986_2605_buf_ack_1, ack => convolve_CP_6526_elements(85)); -- 
    -- CP-element group 86:  join  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	23 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	26 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	25 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_sample_start_
      -- 
    convolve_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(26);
      gj_convolve_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	23 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	281 
    -- CP-element group 87: 	222 
    -- CP-element group 87: 	226 
    -- CP-element group 87: 	274 
    -- CP-element group 87: 	218 
    -- CP-element group 87: 	243 
    -- CP-element group 87: 	247 
    -- CP-element group 87: 	251 
    -- CP-element group 87: 	238 
    -- CP-element group 87: 	230 
    -- CP-element group 87: 	234 
    -- CP-element group 87: 	91 
    -- CP-element group 87: 	175 
    -- CP-element group 87: 	166 
    -- CP-element group 87: 	170 
    -- CP-element group 87: 	146 
    -- CP-element group 87: 	150 
    -- CP-element group 87: 	154 
    -- CP-element group 87: 	158 
    -- CP-element group 87: 	162 
    -- CP-element group 87: 	142 
    -- CP-element group 87: 	212 
    -- CP-element group 87: 	198 
    -- CP-element group 87: 	179 
    -- CP-element group 87: 	183 
    -- CP-element group 87: 	187 
    -- CP-element group 87: 	191 
    -- CP-element group 87: 	205 
    -- CP-element group 87: 	267 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	27 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_update_start_
      -- 
    convolve_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 29) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_markings: IntegerArray(0 to 29)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_delays: IntegerArray(0 to 29) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 30); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(281) & convolve_CP_6526_elements(222) & convolve_CP_6526_elements(226) & convolve_CP_6526_elements(274) & convolve_CP_6526_elements(218) & convolve_CP_6526_elements(243) & convolve_CP_6526_elements(247) & convolve_CP_6526_elements(251) & convolve_CP_6526_elements(238) & convolve_CP_6526_elements(230) & convolve_CP_6526_elements(234) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(175) & convolve_CP_6526_elements(166) & convolve_CP_6526_elements(170) & convolve_CP_6526_elements(146) & convolve_CP_6526_elements(150) & convolve_CP_6526_elements(154) & convolve_CP_6526_elements(158) & convolve_CP_6526_elements(162) & convolve_CP_6526_elements(142) & convolve_CP_6526_elements(212) & convolve_CP_6526_elements(198) & convolve_CP_6526_elements(179) & convolve_CP_6526_elements(183) & convolve_CP_6526_elements(187) & convolve_CP_6526_elements(191) & convolve_CP_6526_elements(205) & convolve_CP_6526_elements(267);
      gj_convolve_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 30, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	25 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_sample_start__ps
      -- 
    convolve_CP_6526_elements(88) <= convolve_CP_6526_elements(25);
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	26 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_sample_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(89) is bound as output of CP function.
    -- CP-element group 90:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	27 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_update_start__ps
      -- 
    convolve_CP_6526_elements(90) <= convolve_CP_6526_elements(27);
    -- CP-element group 91:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	222 
    -- CP-element group 91: 	226 
    -- CP-element group 91: 	272 
    -- CP-element group 91: 	279 
    -- CP-element group 91: 	218 
    -- CP-element group 91: 	245 
    -- CP-element group 91: 	249 
    -- CP-element group 91: 	238 
    -- CP-element group 91: 	241 
    -- CP-element group 91: 	230 
    -- CP-element group 91: 	234 
    -- CP-element group 91: 	24 
    -- CP-element group 91: 	28 
    -- CP-element group 91: 	173 
    -- CP-element group 91: 	177 
    -- CP-element group 91: 	166 
    -- CP-element group 91: 	170 
    -- CP-element group 91: 	146 
    -- CP-element group 91: 	150 
    -- CP-element group 91: 	154 
    -- CP-element group 91: 	158 
    -- CP-element group 91: 	162 
    -- CP-element group 91: 	142 
    -- CP-element group 91: 	210 
    -- CP-element group 91: 	203 
    -- CP-element group 91: 	196 
    -- CP-element group 91: 	181 
    -- CP-element group 91: 	185 
    -- CP-element group 91: 	189 
    -- CP-element group 91: 	265 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	87 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_update_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(91) is bound as output of CP function.
    -- CP-element group 92:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	21 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_loopback_trigger
      -- 
    convolve_CP_6526_elements(92) <= convolve_CP_6526_elements(21);
    -- CP-element group 93:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_loopback_sample_req_ps
      -- CP-element group 93: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_loopback_sample_req
      -- 
    phi_stmt_2606_loopback_sample_req_6791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2606_loopback_sample_req_6791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(93), ack => phi_stmt_2606_req_1); -- 
    -- Element group convolve_CP_6526_elements(93) is bound as output of CP function.
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	22 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_entry_trigger
      -- 
    convolve_CP_6526_elements(94) <= convolve_CP_6526_elements(22);
    -- CP-element group 95:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_entry_sample_req
      -- CP-element group 95: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_entry_sample_req_ps
      -- 
    phi_stmt_2606_entry_sample_req_6794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2606_entry_sample_req_6794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(95), ack => phi_stmt_2606_req_0); -- 
    -- Element group convolve_CP_6526_elements(95) is bound as output of CP function.
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_phi_mux_ack
      -- CP-element group 96: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2606_phi_mux_ack_ps
      -- 
    phi_stmt_2606_phi_mux_ack_6797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2606_ack_0, ack => convolve_CP_6526_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2609_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2609_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2609_sample_start__ps
      -- CP-element group 97: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2609_sample_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(97) is bound as output of CP function.
    -- CP-element group 98:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2609_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2609_update_start__ps
      -- 
    -- Element group convolve_CP_6526_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2609_update_completed__ps
      -- 
    convolve_CP_6526_elements(99) <= convolve_CP_6526_elements(100);
    -- CP-element group 100:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	99 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2609_update_completed_
      -- 
    -- Element group convolve_CP_6526_elements(100) is a control-delay.
    cp_element_100_delay: control_delay_element  generic map(name => " 100_delay", delay_value => 1)  port map(req => convolve_CP_6526_elements(98), ack => convolve_CP_6526_elements(100), clk => clk, reset =>reset);
    -- CP-element group 101:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_sample_start__ps
      -- CP-element group 101: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_Sample/req
      -- CP-element group 101: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_sample_start_
      -- 
    req_6818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(101), ack => n_col_2978_2610_buf_req_0); -- 
    -- Element group convolve_CP_6526_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_update_start_
      -- CP-element group 102: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_Update/req
      -- CP-element group 102: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_update_start__ps
      -- CP-element group 102: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_Update/$entry
      -- 
    req_6823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(102), ack => n_col_2978_2610_buf_req_1); -- 
    -- Element group convolve_CP_6526_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_Sample/ack
      -- CP-element group 103: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_sample_completed__ps
      -- CP-element group 103: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_sample_completed_
      -- 
    ack_6819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_2978_2610_buf_ack_0, ack => convolve_CP_6526_elements(103)); -- 
    -- CP-element group 104:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_update_completed__ps
      -- CP-element group 104: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_col_2610_update_completed_
      -- 
    ack_6824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_2978_2610_buf_ack_1, ack => convolve_CP_6526_elements(104)); -- 
    -- CP-element group 105:  join  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	23 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	26 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	25 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_sample_start_
      -- 
    convolve_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(26);
      gj_convolve_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	23 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: 	288 
    -- CP-element group 106: 	292 
    -- CP-element group 106: 	296 
    -- CP-element group 106: 	175 
    -- CP-element group 106: 	166 
    -- CP-element group 106: 	170 
    -- CP-element group 106: 	307 
    -- CP-element group 106: 	146 
    -- CP-element group 106: 	150 
    -- CP-element group 106: 	154 
    -- CP-element group 106: 	158 
    -- CP-element group 106: 	162 
    -- CP-element group 106: 	142 
    -- CP-element group 106: 	212 
    -- CP-element group 106: 	198 
    -- CP-element group 106: 	179 
    -- CP-element group 106: 	183 
    -- CP-element group 106: 	187 
    -- CP-element group 106: 	191 
    -- CP-element group 106: 	205 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	27 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_update_start_
      -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(108) & convolve_CP_6526_elements(288) & convolve_CP_6526_elements(292) & convolve_CP_6526_elements(296) & convolve_CP_6526_elements(175) & convolve_CP_6526_elements(166) & convolve_CP_6526_elements(170) & convolve_CP_6526_elements(307) & convolve_CP_6526_elements(146) & convolve_CP_6526_elements(150) & convolve_CP_6526_elements(154) & convolve_CP_6526_elements(158) & convolve_CP_6526_elements(162) & convolve_CP_6526_elements(142) & convolve_CP_6526_elements(212) & convolve_CP_6526_elements(198) & convolve_CP_6526_elements(179) & convolve_CP_6526_elements(183) & convolve_CP_6526_elements(187) & convolve_CP_6526_elements(191) & convolve_CP_6526_elements(205);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  join  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	26 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_sample_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(107) is bound as output of CP function.
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	286 
    -- CP-element group 108: 	290 
    -- CP-element group 108: 	294 
    -- CP-element group 108: 	24 
    -- CP-element group 108: 	28 
    -- CP-element group 108: 	173 
    -- CP-element group 108: 	177 
    -- CP-element group 108: 	166 
    -- CP-element group 108: 	170 
    -- CP-element group 108: 	305 
    -- CP-element group 108: 	146 
    -- CP-element group 108: 	150 
    -- CP-element group 108: 	154 
    -- CP-element group 108: 	158 
    -- CP-element group 108: 	162 
    -- CP-element group 108: 	142 
    -- CP-element group 108: 	210 
    -- CP-element group 108: 	203 
    -- CP-element group 108: 	196 
    -- CP-element group 108: 	181 
    -- CP-element group 108: 	185 
    -- CP-element group 108: 	189 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_update_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(108) is bound as output of CP function.
    -- CP-element group 109:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	21 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_loopback_trigger
      -- 
    convolve_CP_6526_elements(109) <= convolve_CP_6526_elements(21);
    -- CP-element group 110:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_loopback_sample_req
      -- CP-element group 110: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_loopback_sample_req_ps
      -- 
    phi_stmt_2611_loopback_sample_req_6835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2611_loopback_sample_req_6835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(110), ack => phi_stmt_2611_req_1); -- 
    -- Element group convolve_CP_6526_elements(110) is bound as output of CP function.
    -- CP-element group 111:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	22 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_entry_trigger
      -- 
    convolve_CP_6526_elements(111) <= convolve_CP_6526_elements(22);
    -- CP-element group 112:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_entry_sample_req
      -- CP-element group 112: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_entry_sample_req_ps
      -- 
    phi_stmt_2611_entry_sample_req_6838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2611_entry_sample_req_6838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(112), ack => phi_stmt_2611_req_0); -- 
    -- Element group convolve_CP_6526_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_phi_mux_ack
      -- CP-element group 113: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2611_phi_mux_ack_ps
      -- 
    phi_stmt_2611_phi_mux_ack_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2611_ack_0, ack => convolve_CP_6526_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2615_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2615_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2615_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2615_sample_completed_
      -- 
    -- Element group convolve_CP_6526_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2615_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2615_update_start_
      -- 
    -- Element group convolve_CP_6526_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2615_update_completed__ps
      -- 
    convolve_CP_6526_elements(116) <= convolve_CP_6526_elements(117);
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2615_update_completed_
      -- 
    -- Element group convolve_CP_6526_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => convolve_CP_6526_elements(115), ack => convolve_CP_6526_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_sample_start__ps
      -- CP-element group 118: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_Sample/req
      -- 
    req_6862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(118), ack => n_num_2967_2616_buf_req_0); -- 
    -- Element group convolve_CP_6526_elements(118) is bound as output of CP function.
    -- CP-element group 119:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_update_start__ps
      -- CP-element group 119: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_update_start_
      -- CP-element group 119: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_Update/req
      -- 
    req_6867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(119), ack => n_num_2967_2616_buf_req_1); -- 
    -- Element group convolve_CP_6526_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (4) 
      -- CP-element group 120: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_sample_completed__ps
      -- CP-element group 120: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_Sample/ack
      -- 
    ack_6863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_2967_2616_buf_ack_0, ack => convolve_CP_6526_elements(120)); -- 
    -- CP-element group 121:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_num_2616_Update/ack
      -- 
    ack_6868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_2967_2616_buf_ack_1, ack => convolve_CP_6526_elements(121)); -- 
    -- CP-element group 122:  join  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	23 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	26 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	25 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_sample_start_
      -- 
    convolve_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(26);
      gj_convolve_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	23 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	288 
    -- CP-element group 123: 	292 
    -- CP-element group 123: 	296 
    -- CP-element group 123: 	127 
    -- CP-element group 123: 	307 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	27 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_update_start_
      -- 
    convolve_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(288) & convolve_CP_6526_elements(292) & convolve_CP_6526_elements(296) & convolve_CP_6526_elements(127) & convolve_CP_6526_elements(307);
      gj_convolve_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	25 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_sample_start__ps
      -- 
    convolve_CP_6526_elements(124) <= convolve_CP_6526_elements(25);
    -- CP-element group 125:  join  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	26 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_sample_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	27 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_update_start__ps
      -- 
    convolve_CP_6526_elements(126) <= convolve_CP_6526_elements(27);
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	286 
    -- CP-element group 127: 	290 
    -- CP-element group 127: 	294 
    -- CP-element group 127: 	24 
    -- CP-element group 127: 	28 
    -- CP-element group 127: 	305 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	123 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_update_completed__ps
      -- 
    -- Element group convolve_CP_6526_elements(127) is bound as output of CP function.
    -- CP-element group 128:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	21 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_loopback_trigger
      -- 
    convolve_CP_6526_elements(128) <= convolve_CP_6526_elements(21);
    -- CP-element group 129:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_loopback_sample_req
      -- CP-element group 129: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_loopback_sample_req_ps
      -- 
    phi_stmt_2617_loopback_sample_req_6879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2617_loopback_sample_req_6879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(129), ack => phi_stmt_2617_req_1); -- 
    -- Element group convolve_CP_6526_elements(129) is bound as output of CP function.
    -- CP-element group 130:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	22 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_entry_trigger
      -- 
    convolve_CP_6526_elements(130) <= convolve_CP_6526_elements(22);
    -- CP-element group 131:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_entry_sample_req
      -- CP-element group 131: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_entry_sample_req_ps
      -- 
    phi_stmt_2617_entry_sample_req_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2617_entry_sample_req_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(131), ack => phi_stmt_2617_req_0); -- 
    -- Element group convolve_CP_6526_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_phi_mux_ack
      -- CP-element group 132: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/phi_stmt_2617_phi_mux_ack_ps
      -- 
    phi_stmt_2617_phi_mux_ack_6885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2617_ack_0, ack => convolve_CP_6526_elements(132)); -- 
    -- CP-element group 133:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2620_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2620_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2620_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2620_sample_completed_
      -- 
    -- Element group convolve_CP_6526_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2620_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2620_update_start_
      -- 
    -- Element group convolve_CP_6526_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2620_update_completed__ps
      -- 
    convolve_CP_6526_elements(135) <= convolve_CP_6526_elements(136);
    -- CP-element group 136:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	135 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_2620_update_completed_
      -- 
    -- Element group convolve_CP_6526_elements(136) is a control-delay.
    cp_element_136_delay: control_delay_element  generic map(name => " 136_delay", delay_value => 1)  port map(req => convolve_CP_6526_elements(134), ack => convolve_CP_6526_elements(136), clk => clk, reset =>reset);
    -- CP-element group 137:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_sample_start__ps
      -- CP-element group 137: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_Sample/req
      -- 
    req_6906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(137), ack => n_chl_2956_2621_buf_req_0); -- 
    -- Element group convolve_CP_6526_elements(137) is bound as output of CP function.
    -- CP-element group 138:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_update_start__ps
      -- CP-element group 138: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_update_start_
      -- CP-element group 138: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_Update/req
      -- 
    req_6911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(138), ack => n_chl_2956_2621_buf_req_1); -- 
    -- Element group convolve_CP_6526_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_sample_completed__ps
      -- CP-element group 139: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_Sample/ack
      -- 
    ack_6907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_2956_2621_buf_ack_0, ack => convolve_CP_6526_elements(139)); -- 
    -- CP-element group 140:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_update_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/R_n_chl_2621_Update/ack
      -- 
    ack_6912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_2956_2621_buf_ack_1, ack => convolve_CP_6526_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	23 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	144 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_Sample/rr
      -- 
    rr_6921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(141), ack => RPIPE_input_pipe1_2634_inst_req_0); -- 
    convolve_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(144);
      gj_convolve_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	108 
    -- CP-element group 142: 	26 
    -- CP-element group 142: 	91 
    -- CP-element group 142: 	143 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	300 
    -- CP-element group 142: 	194 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	106 
    -- CP-element group 142: 	87 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_update_start_
      -- CP-element group 142: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_Update/cr
      -- 
    cr_6926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(142), ack => RPIPE_input_pipe1_2634_inst_req_1); -- 
    convolve_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(143) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(194);
      gj_convolve_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_Sample/ra
      -- 
    ra_6922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_2634_inst_ack_0, ack => convolve_CP_6526_elements(143)); -- 
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	298 
    -- CP-element group 144: 	193 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	29 
    -- CP-element group 144: 	141 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe1_2634_Update/ca
      -- 
    ca_6927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_2634_inst_ack_1, ack => convolve_CP_6526_elements(144)); -- 
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	23 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	148 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_Sample/rr
      -- 
    rr_6935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(145), ack => RPIPE_input_pipe2_2638_inst_req_0); -- 
    convolve_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(148);
      gj_convolve_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	108 
    -- CP-element group 146: 	26 
    -- CP-element group 146: 	91 
    -- CP-element group 146: 	147 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	311 
    -- CP-element group 146: 	300 
    -- CP-element group 146: 	201 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	106 
    -- CP-element group 146: 	87 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_update_start_
      -- CP-element group 146: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_Update/cr
      -- 
    cr_6940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(146), ack => RPIPE_input_pipe2_2638_inst_req_1); -- 
    convolve_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(147) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(201);
      gj_convolve_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_Sample/ra
      -- 
    ra_6936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_2638_inst_ack_0, ack => convolve_CP_6526_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	298 
    -- CP-element group 148: 	309 
    -- CP-element group 148: 	200 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	29 
    -- CP-element group 148: 	48 
    -- CP-element group 148: 	145 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe2_2638_Update/ca
      -- 
    ca_6941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_2638_inst_ack_1, ack => convolve_CP_6526_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	23 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	152 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_Sample/rr
      -- 
    rr_6949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(149), ack => RPIPE_input_pipe3_2642_inst_req_0); -- 
    convolve_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(152);
      gj_convolve_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	108 
    -- CP-element group 150: 	26 
    -- CP-element group 150: 	91 
    -- CP-element group 150: 	151 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	311 
    -- CP-element group 150: 	300 
    -- CP-element group 150: 	208 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	106 
    -- CP-element group 150: 	87 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_update_start_
      -- CP-element group 150: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_Update/cr
      -- 
    cr_6954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(150), ack => RPIPE_input_pipe3_2642_inst_req_1); -- 
    convolve_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(151) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(208);
      gj_convolve_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	150 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_Sample/ra
      -- 
    ra_6950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_2642_inst_ack_0, ack => convolve_CP_6526_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	298 
    -- CP-element group 152: 	309 
    -- CP-element group 152: 	207 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	29 
    -- CP-element group 152: 	48 
    -- CP-element group 152: 	149 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe3_2642_Update/ca
      -- 
    ca_6955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_2642_inst_ack_1, ack => convolve_CP_6526_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	23 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	156 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_Sample/rr
      -- 
    rr_6963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(153), ack => RPIPE_input_pipe4_2646_inst_req_0); -- 
    convolve_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(156);
      gj_convolve_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	108 
    -- CP-element group 154: 	26 
    -- CP-element group 154: 	91 
    -- CP-element group 154: 	155 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	215 
    -- CP-element group 154: 	311 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	106 
    -- CP-element group 154: 	87 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_update_start_
      -- CP-element group 154: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_Update/cr
      -- 
    cr_6968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(154), ack => RPIPE_input_pipe4_2646_inst_req_1); -- 
    convolve_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(155) & convolve_CP_6526_elements(215) & convolve_CP_6526_elements(311);
      gj_convolve_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	154 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_Sample/ra
      -- 
    ra_6964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe4_2646_inst_ack_0, ack => convolve_CP_6526_elements(155)); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	309 
    -- CP-element group 156: 	214 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	48 
    -- CP-element group 156: 	153 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_input_pipe4_2646_Update/ca
      -- 
    ca_6969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe4_2646_inst_ack_1, ack => convolve_CP_6526_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	23 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	160 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_Sample/rr
      -- 
    rr_6977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(157), ack => RPIPE_xxconvolvexxconv_ip1_2650_inst_req_0); -- 
    convolve_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(160);
      gj_convolve_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	108 
    -- CP-element group 158: 	26 
    -- CP-element group 158: 	91 
    -- CP-element group 158: 	159 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	300 
    -- CP-element group 158: 	194 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	106 
    -- CP-element group 158: 	87 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_update_start_
      -- CP-element group 158: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_Update/cr
      -- 
    cr_6982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(158), ack => RPIPE_xxconvolvexxconv_ip1_2650_inst_req_1); -- 
    convolve_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(159) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(194);
      gj_convolve_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	158 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_Sample/ra
      -- 
    ra_6978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_2650_inst_ack_0, ack => convolve_CP_6526_elements(159)); -- 
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	298 
    -- CP-element group 160: 	193 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	29 
    -- CP-element group 160: 	157 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip1_2650_Update/ca
      -- 
    ca_6983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_2650_inst_ack_1, ack => convolve_CP_6526_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	23 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	164 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_Sample/rr
      -- 
    rr_6991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(161), ack => RPIPE_xxconvolvexxconv_ip2_2654_inst_req_0); -- 
    convolve_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(164);
      gj_convolve_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	108 
    -- CP-element group 162: 	26 
    -- CP-element group 162: 	91 
    -- CP-element group 162: 	163 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	311 
    -- CP-element group 162: 	300 
    -- CP-element group 162: 	201 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	106 
    -- CP-element group 162: 	87 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_update_start_
      -- CP-element group 162: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_Update/cr
      -- 
    cr_6996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(162), ack => RPIPE_xxconvolvexxconv_ip2_2654_inst_req_1); -- 
    convolve_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(163) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(201);
      gj_convolve_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	162 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_Sample/ra
      -- 
    ra_6992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_2654_inst_ack_0, ack => convolve_CP_6526_elements(163)); -- 
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	298 
    -- CP-element group 164: 	309 
    -- CP-element group 164: 	200 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	29 
    -- CP-element group 164: 	48 
    -- CP-element group 164: 	161 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip2_2654_Update/ca
      -- 
    ca_6997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_2654_inst_ack_1, ack => convolve_CP_6526_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	23 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	168 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_Sample/rr
      -- 
    rr_7005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(165), ack => RPIPE_xxconvolvexxconv_ip3_2658_inst_req_0); -- 
    convolve_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(168);
      gj_convolve_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	108 
    -- CP-element group 166: 	26 
    -- CP-element group 166: 	91 
    -- CP-element group 166: 	167 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	311 
    -- CP-element group 166: 	300 
    -- CP-element group 166: 	208 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	106 
    -- CP-element group 166: 	87 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_update_start_
      -- CP-element group 166: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_Update/cr
      -- 
    cr_7010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(166), ack => RPIPE_xxconvolvexxconv_ip3_2658_inst_req_1); -- 
    convolve_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(167) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(208);
      gj_convolve_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	166 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_Sample/ra
      -- 
    ra_7006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_2658_inst_ack_0, ack => convolve_CP_6526_elements(167)); -- 
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	298 
    -- CP-element group 168: 	309 
    -- CP-element group 168: 	207 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	29 
    -- CP-element group 168: 	48 
    -- CP-element group 168: 	165 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip3_2658_Update/ca
      -- 
    ca_7011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_2658_inst_ack_1, ack => convolve_CP_6526_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	23 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	172 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_Sample/rr
      -- 
    rr_7019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(169), ack => RPIPE_xxconvolvexxconv_ip4_2662_inst_req_0); -- 
    convolve_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(172);
      gj_convolve_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	108 
    -- CP-element group 170: 	26 
    -- CP-element group 170: 	91 
    -- CP-element group 170: 	171 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	215 
    -- CP-element group 170: 	311 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	106 
    -- CP-element group 170: 	87 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_update_start_
      -- CP-element group 170: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_Update/cr
      -- 
    cr_7024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(170), ack => RPIPE_xxconvolvexxconv_ip4_2662_inst_req_1); -- 
    convolve_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(171) & convolve_CP_6526_elements(215) & convolve_CP_6526_elements(311);
      gj_convolve_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	170 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_Sample/ra
      -- 
    ra_7020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip4_2662_inst_ack_0, ack => convolve_CP_6526_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	309 
    -- CP-element group 172: 	214 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	48 
    -- CP-element group 172: 	169 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_ip4_2662_Update/ca
      -- 
    ca_7025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip4_2662_inst_ack_1, ack => convolve_CP_6526_elements(172)); -- 
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	108 
    -- CP-element group 173: 	91 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_Sample/req
      -- 
    req_7033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(173), ack => W_read_ip_2608_delayed_1_0_2664_inst_req_0); -- 
    convolve_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(175);
      gj_convolve_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	26 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: 	300 
    -- CP-element group 174: 	194 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_update_start_
      -- CP-element group 174: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_Update/req
      -- 
    req_7038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(174), ack => W_read_ip_2608_delayed_1_0_2664_inst_req_1); -- 
    convolve_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(176) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(194);
      gj_convolve_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	106 
    -- CP-element group 175: 	87 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_Sample/ack
      -- 
    ack_7034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2608_delayed_1_0_2664_inst_ack_0, ack => convolve_CP_6526_elements(175)); -- 
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	298 
    -- CP-element group 176: 	193 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	29 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2666_Update/ack
      -- 
    ack_7039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2608_delayed_1_0_2664_inst_ack_1, ack => convolve_CP_6526_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	108 
    -- CP-element group 177: 	91 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_Sample/req
      -- 
    req_7047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(177), ack => W_read_ip_2614_delayed_1_0_2673_inst_req_0); -- 
    convolve_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(179);
      gj_convolve_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	26 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	311 
    -- CP-element group 178: 	300 
    -- CP-element group 178: 	201 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_update_start_
      -- CP-element group 178: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_Update/req
      -- 
    req_7052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(178), ack => W_read_ip_2614_delayed_1_0_2673_inst_req_1); -- 
    convolve_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(201) & convolve_CP_6526_elements(180);
      gj_convolve_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	106 
    -- CP-element group 179: 	87 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_Sample/ack
      -- 
    ack_7048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2614_delayed_1_0_2673_inst_ack_0, ack => convolve_CP_6526_elements(179)); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	298 
    -- CP-element group 180: 	309 
    -- CP-element group 180: 	200 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	29 
    -- CP-element group 180: 	48 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2675_Update/ack
      -- 
    ack_7053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2614_delayed_1_0_2673_inst_ack_1, ack => convolve_CP_6526_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	108 
    -- CP-element group 181: 	91 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_Sample/req
      -- 
    req_7061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(181), ack => W_read_ip_2620_delayed_1_0_2682_inst_req_0); -- 
    convolve_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(183);
      gj_convolve_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	26 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	311 
    -- CP-element group 182: 	300 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	208 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_update_start_
      -- CP-element group 182: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_Update/req
      -- 
    req_7066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(182), ack => W_read_ip_2620_delayed_1_0_2682_inst_req_1); -- 
    convolve_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(184) & convolve_CP_6526_elements(208);
      gj_convolve_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	106 
    -- CP-element group 183: 	87 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_Sample/ack
      -- 
    ack_7062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2620_delayed_1_0_2682_inst_ack_0, ack => convolve_CP_6526_elements(183)); -- 
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	298 
    -- CP-element group 184: 	309 
    -- CP-element group 184: 	207 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	29 
    -- CP-element group 184: 	48 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2684_Update/ack
      -- 
    ack_7067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2620_delayed_1_0_2682_inst_ack_1, ack => convolve_CP_6526_elements(184)); -- 
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	108 
    -- CP-element group 185: 	91 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_Sample/req
      -- 
    req_7075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(185), ack => W_read_ip_2626_delayed_1_0_2691_inst_req_0); -- 
    convolve_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(187);
      gj_convolve_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	26 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	215 
    -- CP-element group 186: 	311 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_update_start_
      -- CP-element group 186: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_Update/req
      -- 
    req_7080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(186), ack => W_read_ip_2626_delayed_1_0_2691_inst_req_1); -- 
    convolve_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(215) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(188);
      gj_convolve_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	106 
    -- CP-element group 187: 	87 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_Sample/ack
      -- 
    ack_7076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2626_delayed_1_0_2691_inst_ack_0, ack => convolve_CP_6526_elements(187)); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	309 
    -- CP-element group 188: 	214 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	48 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2693_Update/ack
      -- 
    ack_7081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_2626_delayed_1_0_2691_inst_ack_1, ack => convolve_CP_6526_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	108 
    -- CP-element group 189: 	91 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_Sample/req
      -- 
    req_7089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(189), ack => W_write_input_2640_delayed_1_0_2709_inst_req_0); -- 
    convolve_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(191);
      gj_convolve_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_update_start_
      -- CP-element group 190: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_Update/req
      -- 
    req_7094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(190), ack => W_write_input_2640_delayed_1_0_2709_inst_req_1); -- 
    convolve_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(192) & convolve_CP_6526_elements(194);
      gj_convolve_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	106 
    -- CP-element group 191: 	87 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_Sample/ack
      -- 
    ack_7090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2640_delayed_1_0_2709_inst_ack_0, ack => convolve_CP_6526_elements(191)); -- 
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2711_Update/ack
      -- 
    ack_7095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2640_delayed_1_0_2709_inst_ack_1, ack => convolve_CP_6526_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	176 
    -- CP-element group 193: 	160 
    -- CP-element group 193: 	144 
    -- CP-element group 193: 	192 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_Sample/req
      -- 
    req_7103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(193), ack => WPIPE_xxconvolvexxconv_ip1_2713_inst_req_0); -- 
    convolve_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(176) & convolve_CP_6526_elements(160) & convolve_CP_6526_elements(144) & convolve_CP_6526_elements(192) & convolve_CP_6526_elements(195);
      gj_convolve_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	174 
    -- CP-element group 194: 	158 
    -- CP-element group 194: 	142 
    -- CP-element group 194: 	190 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_update_start_
      -- CP-element group 194: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_Update/req
      -- 
    ack_7104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2713_inst_ack_0, ack => convolve_CP_6526_elements(194)); -- 
    req_7108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(194), ack => WPIPE_xxconvolvexxconv_ip1_2713_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	317 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip1_2713_Update/ack
      -- 
    ack_7109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2713_inst_ack_1, ack => convolve_CP_6526_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	108 
    -- CP-element group 196: 	91 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_Sample/req
      -- 
    req_7117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(196), ack => W_write_input_2644_delayed_1_0_2716_inst_req_0); -- 
    convolve_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(198);
      gj_convolve_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_update_start_
      -- CP-element group 197: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_Update/req
      -- 
    req_7122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(197), ack => W_write_input_2644_delayed_1_0_2716_inst_req_1); -- 
    convolve_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(199) & convolve_CP_6526_elements(201);
      gj_convolve_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	106 
    -- CP-element group 198: 	87 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_Sample/ack
      -- 
    ack_7118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2644_delayed_1_0_2716_inst_ack_0, ack => convolve_CP_6526_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2718_Update/ack
      -- 
    ack_7123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2644_delayed_1_0_2716_inst_ack_1, ack => convolve_CP_6526_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	148 
    -- CP-element group 200: 	164 
    -- CP-element group 200: 	199 
    -- CP-element group 200: 	180 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_Sample/req
      -- 
    req_7131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(200), ack => WPIPE_xxconvolvexxconv_ip2_2720_inst_req_0); -- 
    convolve_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(148) & convolve_CP_6526_elements(164) & convolve_CP_6526_elements(199) & convolve_CP_6526_elements(180) & convolve_CP_6526_elements(202);
      gj_convolve_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	178 
    -- CP-element group 201: 	146 
    -- CP-element group 201: 	162 
    -- CP-element group 201: 	197 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_Update/req
      -- CP-element group 201: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_update_start_
      -- CP-element group 201: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_Sample/ack
      -- 
    ack_7132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2720_inst_ack_0, ack => convolve_CP_6526_elements(201)); -- 
    req_7136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(201), ack => WPIPE_xxconvolvexxconv_ip2_2720_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	317 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_Update/ack
      -- CP-element group 202: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip2_2720_update_completed_
      -- 
    ack_7137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2720_inst_ack_1, ack => convolve_CP_6526_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	108 
    -- CP-element group 203: 	91 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_Sample/req
      -- CP-element group 203: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_sample_start_
      -- 
    req_7145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(203), ack => W_write_input_2648_delayed_1_0_2723_inst_req_0); -- 
    convolve_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(205);
      gj_convolve_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: 	208 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_update_start_
      -- CP-element group 204: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_Update/req
      -- CP-element group 204: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_Update/$entry
      -- 
    req_7150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(204), ack => W_write_input_2648_delayed_1_0_2723_inst_req_1); -- 
    convolve_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(206) & convolve_CP_6526_elements(208);
      gj_convolve_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	106 
    -- CP-element group 205: 	87 
    -- CP-element group 205: 	203 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_Sample/ack
      -- 
    ack_7146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2648_delayed_1_0_2723_inst_ack_0, ack => convolve_CP_6526_elements(205)); -- 
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_Update/ack
      -- CP-element group 206: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2725_Update/$exit
      -- 
    ack_7151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2648_delayed_1_0_2723_inst_ack_1, ack => convolve_CP_6526_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	168 
    -- CP-element group 207: 	152 
    -- CP-element group 207: 	184 
    -- CP-element group 207: 	206 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_Sample/req
      -- 
    req_7159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(207), ack => WPIPE_xxconvolvexxconv_ip3_2727_inst_req_0); -- 
    convolve_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(168) & convolve_CP_6526_elements(152) & convolve_CP_6526_elements(184) & convolve_CP_6526_elements(206) & convolve_CP_6526_elements(209);
      gj_convolve_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	166 
    -- CP-element group 208: 	150 
    -- CP-element group 208: 	182 
    -- CP-element group 208: 	204 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_update_start_
      -- CP-element group 208: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_Update/req
      -- CP-element group 208: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_Sample/ack
      -- CP-element group 208: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_Sample/$exit
      -- 
    ack_7160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2727_inst_ack_0, ack => convolve_CP_6526_elements(208)); -- 
    req_7164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(208), ack => WPIPE_xxconvolvexxconv_ip3_2727_inst_req_1); -- 
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	317 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_Update/ack
      -- CP-element group 209: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip3_2727_Update/$exit
      -- 
    ack_7165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2727_inst_ack_1, ack => convolve_CP_6526_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	108 
    -- CP-element group 210: 	91 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_Sample/req
      -- CP-element group 210: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_sample_start_
      -- 
    req_7173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(210), ack => W_write_input_2652_delayed_1_0_2730_inst_req_0); -- 
    convolve_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(212);
      gj_convolve_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	215 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_Update/req
      -- CP-element group 211: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_update_start_
      -- 
    req_7178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(211), ack => W_write_input_2652_delayed_1_0_2730_inst_req_1); -- 
    convolve_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(215) & convolve_CP_6526_elements(213);
      gj_convolve_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	106 
    -- CP-element group 212: 	87 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_Sample/ack
      -- CP-element group 212: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_sample_completed_
      -- 
    ack_7174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2652_delayed_1_0_2730_inst_ack_0, ack => convolve_CP_6526_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_Update/ack
      -- CP-element group 213: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2732_update_completed_
      -- 
    ack_7179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_2652_delayed_1_0_2730_inst_ack_1, ack => convolve_CP_6526_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	172 
    -- CP-element group 214: 	156 
    -- CP-element group 214: 	213 
    -- CP-element group 214: 	188 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_Sample/req
      -- CP-element group 214: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_Sample/$entry
      -- 
    req_7187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(214), ack => WPIPE_xxconvolvexxconv_ip4_2734_inst_req_0); -- 
    convolve_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(172) & convolve_CP_6526_elements(156) & convolve_CP_6526_elements(213) & convolve_CP_6526_elements(188) & convolve_CP_6526_elements(216);
      gj_convolve_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	170 
    -- CP-element group 215: 	154 
    -- CP-element group 215: 	211 
    -- CP-element group 215: 	186 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_update_start_
      -- CP-element group 215: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_Update/req
      -- CP-element group 215: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_Update/$entry
      -- 
    ack_7188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip4_2734_inst_ack_0, ack => convolve_CP_6526_elements(215)); -- 
    req_7192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(215), ack => WPIPE_xxconvolvexxconv_ip4_2734_inst_req_1); -- 
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	317 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_Update/ack
      -- CP-element group 216: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_ip4_2734_Update/$exit
      -- 
    ack_7193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip4_2734_inst_ack_1, ack => convolve_CP_6526_elements(216)); -- 
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	23 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	220 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_Sample/rr
      -- CP-element group 217: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_Sample/$entry
      -- CP-element group 217: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_sample_start_
      -- 
    rr_7201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(217), ack => RPIPE_kernel_pipe1_2764_inst_req_0); -- 
    convolve_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(220);
      gj_convolve_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	219 
    -- CP-element group 218: 	26 
    -- CP-element group 218: 	72 
    -- CP-element group 218: 	91 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	270 
    -- CP-element group 218: 	311 
    -- CP-element group 218: 	300 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	68 
    -- CP-element group 218: 	87 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_update_start_
      -- 
    cr_7206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(218), ack => RPIPE_kernel_pipe1_2764_inst_req_1); -- 
    convolve_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(219) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(270) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	218 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_Sample/ra
      -- CP-element group 219: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_sample_completed_
      -- 
    ra_7202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2764_inst_ack_0, ack => convolve_CP_6526_elements(219)); -- 
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	269 
    -- CP-element group 220: 	298 
    -- CP-element group 220: 	309 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	217 
    -- CP-element group 220: 	29 
    -- CP-element group 220: 	48 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_Update/ca
      -- CP-element group 220: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe1_2764_Update/$exit
      -- 
    ca_7207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2764_inst_ack_1, ack => convolve_CP_6526_elements(220)); -- 
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	23 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	224 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_Sample/rr
      -- CP-element group 221: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_sample_start_
      -- 
    rr_7215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(221), ack => RPIPE_kernel_pipe2_2768_inst_req_0); -- 
    convolve_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(224);
      gj_convolve_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	223 
    -- CP-element group 222: 	26 
    -- CP-element group 222: 	72 
    -- CP-element group 222: 	91 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	277 
    -- CP-element group 222: 	311 
    -- CP-element group 222: 	300 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	68 
    -- CP-element group 222: 	87 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_Update/cr
      -- CP-element group 222: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_Update/$entry
      -- CP-element group 222: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_update_start_
      -- 
    cr_7220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(222), ack => RPIPE_kernel_pipe2_2768_inst_req_1); -- 
    convolve_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(223) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(277) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	222 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_Sample/ra
      -- CP-element group 223: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_sample_completed_
      -- 
    ra_7216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2768_inst_ack_0, ack => convolve_CP_6526_elements(223)); -- 
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	276 
    -- CP-element group 224: 	298 
    -- CP-element group 224: 	309 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	221 
    -- CP-element group 224: 	29 
    -- CP-element group 224: 	48 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_Update/ca
      -- CP-element group 224: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe2_2768_update_completed_
      -- 
    ca_7221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2768_inst_ack_1, ack => convolve_CP_6526_elements(224)); -- 
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	23 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	228 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_Sample/rr
      -- 
    rr_7229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(225), ack => RPIPE_kernel_pipe3_2772_inst_req_0); -- 
    convolve_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(228);
      gj_convolve_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	227 
    -- CP-element group 226: 	26 
    -- CP-element group 226: 	72 
    -- CP-element group 226: 	91 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	284 
    -- CP-element group 226: 	311 
    -- CP-element group 226: 	300 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	68 
    -- CP-element group 226: 	87 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_update_start_
      -- CP-element group 226: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_Update/cr
      -- 
    cr_7234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(226), ack => RPIPE_kernel_pipe3_2772_inst_req_1); -- 
    convolve_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(227) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(284) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	226 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_Sample/ra
      -- 
    ra_7230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2772_inst_ack_0, ack => convolve_CP_6526_elements(227)); -- 
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	283 
    -- CP-element group 228: 	298 
    -- CP-element group 228: 	309 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	225 
    -- CP-element group 228: 	29 
    -- CP-element group 228: 	48 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_kernel_pipe3_2772_Update/ca
      -- 
    ca_7235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2772_inst_ack_1, ack => convolve_CP_6526_elements(228)); -- 
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	23 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	232 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_Sample/rr
      -- CP-element group 229: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_sample_start_
      -- 
    rr_7243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(229), ack => RPIPE_xxconvolvexxconv_k1_2776_inst_req_0); -- 
    convolve_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(232);
      gj_convolve_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	231 
    -- CP-element group 230: 	26 
    -- CP-element group 230: 	72 
    -- CP-element group 230: 	91 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	270 
    -- CP-element group 230: 	311 
    -- CP-element group 230: 	300 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	68 
    -- CP-element group 230: 	87 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_Update/cr
      -- CP-element group 230: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_update_start_
      -- 
    cr_7248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(230), ack => RPIPE_xxconvolvexxconv_k1_2776_inst_req_1); -- 
    convolve_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(231) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(270) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	230 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_Sample/ra
      -- CP-element group 231: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_sample_completed_
      -- 
    ra_7244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2776_inst_ack_0, ack => convolve_CP_6526_elements(231)); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	269 
    -- CP-element group 232: 	298 
    -- CP-element group 232: 	309 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	229 
    -- CP-element group 232: 	29 
    -- CP-element group 232: 	48 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_Update/ca
      -- CP-element group 232: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k1_2776_update_completed_
      -- 
    ca_7249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2776_inst_ack_1, ack => convolve_CP_6526_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	23 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	236 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_Sample/rr
      -- CP-element group 233: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_sample_start_
      -- 
    rr_7257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(233), ack => RPIPE_xxconvolvexxconv_k2_2780_inst_req_0); -- 
    convolve_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(236);
      gj_convolve_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	26 
    -- CP-element group 234: 	72 
    -- CP-element group 234: 	91 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	277 
    -- CP-element group 234: 	311 
    -- CP-element group 234: 	300 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	68 
    -- CP-element group 234: 	87 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_update_start_
      -- 
    cr_7262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(234), ack => RPIPE_xxconvolvexxconv_k2_2780_inst_req_1); -- 
    convolve_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(235) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(277) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	234 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_Sample/ra
      -- CP-element group 235: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_sample_completed_
      -- 
    ra_7258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2780_inst_ack_0, ack => convolve_CP_6526_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	276 
    -- CP-element group 236: 	298 
    -- CP-element group 236: 	309 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	233 
    -- CP-element group 236: 	29 
    -- CP-element group 236: 	48 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_Update/ca
      -- CP-element group 236: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k2_2780_update_completed_
      -- 
    ca_7263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2780_inst_ack_1, ack => convolve_CP_6526_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	23 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	240 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_Sample/rr
      -- CP-element group 237: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_sample_start_
      -- 
    rr_7271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(237), ack => RPIPE_xxconvolvexxconv_k3_2784_inst_req_0); -- 
    convolve_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(240);
      gj_convolve_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: 	26 
    -- CP-element group 238: 	72 
    -- CP-element group 238: 	91 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	284 
    -- CP-element group 238: 	311 
    -- CP-element group 238: 	300 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	68 
    -- CP-element group 238: 	87 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_Update/cr
      -- CP-element group 238: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_update_start_
      -- 
    cr_7276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(238), ack => RPIPE_xxconvolvexxconv_k3_2784_inst_req_1); -- 
    convolve_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 15,2 => 15,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(239) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(284) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	238 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_Sample/ra
      -- CP-element group 239: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_sample_completed_
      -- 
    ra_7272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2784_inst_ack_0, ack => convolve_CP_6526_elements(239)); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	283 
    -- CP-element group 240: 	298 
    -- CP-element group 240: 	309 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	237 
    -- CP-element group 240: 	29 
    -- CP-element group 240: 	48 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_Update/ca
      -- CP-element group 240: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/RPIPE_xxconvolvexxconv_k3_2784_update_completed_
      -- 
    ca_7277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2784_inst_ack_1, ack => convolve_CP_6526_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	72 
    -- CP-element group 241: 	91 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_Sample/req
      -- 
    req_7285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(241), ack => W_read_k_2706_delayed_1_0_2786_inst_req_0); -- 
    convolve_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(243);
      gj_convolve_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	26 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	270 
    -- CP-element group 242: 	244 
    -- CP-element group 242: 	311 
    -- CP-element group 242: 	300 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_update_start_
      -- CP-element group 242: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_Update/req
      -- CP-element group 242: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_Update/$entry
      -- 
    req_7290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(242), ack => W_read_k_2706_delayed_1_0_2786_inst_req_1); -- 
    convolve_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(270) & convolve_CP_6526_elements(244) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: 	68 
    -- CP-element group 243: 	87 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_Sample/ack
      -- 
    ack_7286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2706_delayed_1_0_2786_inst_ack_0, ack => convolve_CP_6526_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	269 
    -- CP-element group 244: 	298 
    -- CP-element group 244: 	309 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	29 
    -- CP-element group 244: 	48 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2788_Update/$exit
      -- 
    ack_7291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2706_delayed_1_0_2786_inst_ack_1, ack => convolve_CP_6526_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	72 
    -- CP-element group 245: 	91 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_Sample/req
      -- CP-element group 245: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_sample_start_
      -- 
    req_7299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(245), ack => W_read_k_2712_delayed_1_0_2795_inst_req_0); -- 
    convolve_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(247);
      gj_convolve_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	26 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	277 
    -- CP-element group 246: 	248 
    -- CP-element group 246: 	311 
    -- CP-element group 246: 	300 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_Update/req
      -- CP-element group 246: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_update_start_
      -- 
    req_7304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(246), ack => W_read_k_2712_delayed_1_0_2795_inst_req_1); -- 
    convolve_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(277) & convolve_CP_6526_elements(248) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: 	68 
    -- CP-element group 247: 	87 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_sample_completed_
      -- 
    ack_7300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2712_delayed_1_0_2795_inst_ack_0, ack => convolve_CP_6526_elements(247)); -- 
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	276 
    -- CP-element group 248: 	298 
    -- CP-element group 248: 	309 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: 	29 
    -- CP-element group 248: 	48 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2797_update_completed_
      -- 
    ack_7305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2712_delayed_1_0_2795_inst_ack_1, ack => convolve_CP_6526_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	72 
    -- CP-element group 249: 	91 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_Sample/req
      -- CP-element group 249: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_sample_start_
      -- 
    req_7313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(249), ack => W_read_k_2718_delayed_1_0_2804_inst_req_0); -- 
    convolve_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(251);
      gj_convolve_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	26 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	284 
    -- CP-element group 250: 	252 
    -- CP-element group 250: 	311 
    -- CP-element group 250: 	300 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_Update/req
      -- CP-element group 250: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_update_start_
      -- 
    req_7318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(250), ack => W_read_k_2718_delayed_1_0_2804_inst_req_1); -- 
    convolve_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(284) & convolve_CP_6526_elements(252) & convolve_CP_6526_elements(311) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: 	68 
    -- CP-element group 251: 	87 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_sample_completed_
      -- 
    ack_7314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2718_delayed_1_0_2804_inst_ack_0, ack => convolve_CP_6526_elements(251)); -- 
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	283 
    -- CP-element group 252: 	298 
    -- CP-element group 252: 	309 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	29 
    -- CP-element group 252: 	48 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2806_update_completed_
      -- 
    ack_7319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2718_delayed_1_0_2804_inst_ack_1, ack => convolve_CP_6526_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	34 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_Sample/req
      -- CP-element group 253: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_Sample/$entry
      -- 
    req_7327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(253), ack => W_acc1_2772_delayed_1_0_2861_inst_req_0); -- 
    convolve_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(34) & convolve_CP_6526_elements(255);
      gj_convolve_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	26 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: 	300 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_update_start_
      -- CP-element group 254: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_Update/req
      -- CP-element group 254: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_Update/$entry
      -- 
    req_7332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(254), ack => W_acc1_2772_delayed_1_0_2861_inst_req_1); -- 
    convolve_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(256) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: 	30 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_Sample/$exit
      -- 
    ack_7328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc1_2772_delayed_1_0_2861_inst_ack_0, ack => convolve_CP_6526_elements(255)); -- 
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	298 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	29 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2863_Update/$exit
      -- 
    ack_7333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc1_2772_delayed_1_0_2861_inst_ack_1, ack => convolve_CP_6526_elements(256)); -- 
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	53 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_Sample/req
      -- CP-element group 257: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_Sample/$entry
      -- CP-element group 257: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_sample_start_
      -- 
    req_7341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(257), ack => W_acc2_2781_delayed_1_0_2873_inst_req_0); -- 
    convolve_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(53) & convolve_CP_6526_elements(259);
      gj_convolve_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	26 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: 	311 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_Update/req
      -- CP-element group 258: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_update_start_
      -- 
    req_7346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(258), ack => W_acc2_2781_delayed_1_0_2873_inst_req_1); -- 
    convolve_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(260) & convolve_CP_6526_elements(311);
      gj_convolve_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: 	49 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_sample_completed_
      -- 
    ack_7342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc2_2781_delayed_1_0_2873_inst_ack_0, ack => convolve_CP_6526_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	309 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	48 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2875_update_completed_
      -- 
    ack_7347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc2_2781_delayed_1_0_2873_inst_ack_1, ack => convolve_CP_6526_elements(260)); -- 
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	23 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_Sample/rr
      -- CP-element group 261: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_Sample/$entry
      -- 
    rr_7355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(261), ack => SUB_u16_u16_2910_inst_req_0); -- 
    convolve_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(23) & convolve_CP_6526_elements(263);
      gj_convolve_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	281 
    -- CP-element group 262: 	274 
    -- CP-element group 262: 	264 
    -- CP-element group 262: 	267 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_update_start_
      -- 
    cr_7360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(262), ack => SUB_u16_u16_2910_inst_req_1); -- 
    convolve_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(281) & convolve_CP_6526_elements(274) & convolve_CP_6526_elements(264) & convolve_CP_6526_elements(267);
      gj_convolve_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_Sample/ra
      -- CP-element group 263: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_sample_completed_
      -- 
    ra_7356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2910_inst_ack_0, ack => convolve_CP_6526_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	272 
    -- CP-element group 264: 	279 
    -- CP-element group 264: 	24 
    -- CP-element group 264: 	265 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_Update/ca
      -- CP-element group 264: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/SUB_u16_u16_2910_update_completed_
      -- 
    ca_7361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2910_inst_ack_1, ack => convolve_CP_6526_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	72 
    -- CP-element group 265: 	91 
    -- CP-element group 265: 	264 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_Sample/req
      -- CP-element group 265: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_sample_start_
      -- 
    req_7369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(265), ack => W_store_kernel_2829_delayed_1_0_2928_inst_req_0); -- 
    convolve_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(264) & convolve_CP_6526_elements(267);
      gj_convolve_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: 	270 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_update_start_
      -- CP-element group 266: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_Update/req
      -- CP-element group 266: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_Update/$entry
      -- 
    req_7374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(266), ack => W_store_kernel_2829_delayed_1_0_2928_inst_req_1); -- 
    convolve_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(268) & convolve_CP_6526_elements(270);
      gj_convolve_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	68 
    -- CP-element group 267: 	87 
    -- CP-element group 267: 	262 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_Sample/ack
      -- 
    ack_7370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2829_delayed_1_0_2928_inst_ack_0, ack => convolve_CP_6526_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2930_Update/$exit
      -- 
    ack_7375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2829_delayed_1_0_2928_inst_ack_1, ack => convolve_CP_6526_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: 	220 
    -- CP-element group 269: 	244 
    -- CP-element group 269: 	232 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_Sample/req
      -- CP-element group 269: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_sample_start_
      -- 
    req_7383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(269), ack => WPIPE_xxconvolvexxconv_k1_2932_inst_req_0); -- 
    convolve_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(268) & convolve_CP_6526_elements(220) & convolve_CP_6526_elements(244) & convolve_CP_6526_elements(232) & convolve_CP_6526_elements(271);
      gj_convolve_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	218 
    -- CP-element group 270: 	242 
    -- CP-element group 270: 	230 
    -- CP-element group 270: 	266 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_Update/req
      -- CP-element group 270: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_Sample/ack
      -- CP-element group 270: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_update_start_
      -- CP-element group 270: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_sample_completed_
      -- 
    ack_7384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_2932_inst_ack_0, ack => convolve_CP_6526_elements(270)); -- 
    req_7388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(270), ack => WPIPE_xxconvolvexxconv_k1_2932_inst_req_1); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	317 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_Update/ack
      -- CP-element group 271: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k1_2932_update_completed_
      -- 
    ack_7389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_2932_inst_ack_1, ack => convolve_CP_6526_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	72 
    -- CP-element group 272: 	91 
    -- CP-element group 272: 	264 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_sample_start_
      -- 
    req_7397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(272), ack => W_store_kernel_2833_delayed_1_0_2935_inst_req_0); -- 
    convolve_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(264) & convolve_CP_6526_elements(274);
      gj_convolve_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: 	277 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_Update/req
      -- CP-element group 273: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_update_start_
      -- 
    req_7402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(273), ack => W_store_kernel_2833_delayed_1_0_2935_inst_req_1); -- 
    convolve_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(275) & convolve_CP_6526_elements(277);
      gj_convolve_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: 	68 
    -- CP-element group 274: 	87 
    -- CP-element group 274: 	262 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_Sample/ack
      -- CP-element group 274: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_sample_completed_
      -- 
    ack_7398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2833_delayed_1_0_2935_inst_ack_0, ack => convolve_CP_6526_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_Update/ack
      -- CP-element group 275: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2937_update_completed_
      -- 
    ack_7403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2833_delayed_1_0_2935_inst_ack_1, ack => convolve_CP_6526_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	224 
    -- CP-element group 276: 	275 
    -- CP-element group 276: 	248 
    -- CP-element group 276: 	236 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_sample_start_
      -- 
    req_7411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(276), ack => WPIPE_xxconvolvexxconv_k2_2939_inst_req_0); -- 
    convolve_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(224) & convolve_CP_6526_elements(275) & convolve_CP_6526_elements(248) & convolve_CP_6526_elements(236) & convolve_CP_6526_elements(278);
      gj_convolve_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	222 
    -- CP-element group 277: 	273 
    -- CP-element group 277: 	246 
    -- CP-element group 277: 	234 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_Update/req
      -- CP-element group 277: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_update_start_
      -- CP-element group 277: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_sample_completed_
      -- 
    ack_7412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_2939_inst_ack_0, ack => convolve_CP_6526_elements(277)); -- 
    req_7416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(277), ack => WPIPE_xxconvolvexxconv_k2_2939_inst_req_1); -- 
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	317 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k2_2939_update_completed_
      -- 
    ack_7417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_2939_inst_ack_1, ack => convolve_CP_6526_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	72 
    -- CP-element group 279: 	91 
    -- CP-element group 279: 	264 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_Sample/req
      -- CP-element group 279: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_sample_start_
      -- 
    req_7425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(279), ack => W_store_kernel_2837_delayed_1_0_2942_inst_req_0); -- 
    convolve_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(72) & convolve_CP_6526_elements(91) & convolve_CP_6526_elements(264) & convolve_CP_6526_elements(281);
      gj_convolve_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	282 
    -- CP-element group 280: 	284 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_Update/req
      -- CP-element group 280: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_Update/$entry
      -- CP-element group 280: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_update_start_
      -- 
    req_7430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(280), ack => W_store_kernel_2837_delayed_1_0_2942_inst_req_1); -- 
    convolve_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(282) & convolve_CP_6526_elements(284);
      gj_convolve_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281: marked-successors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: 	68 
    -- CP-element group 281: 	87 
    -- CP-element group 281: 	262 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_Sample/ack
      -- CP-element group 281: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_sample_completed_
      -- 
    ack_7426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2837_delayed_1_0_2942_inst_ack_0, ack => convolve_CP_6526_elements(281)); -- 
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2944_Update/ack
      -- 
    ack_7431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2837_delayed_1_0_2942_inst_ack_1, ack => convolve_CP_6526_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: 	252 
    -- CP-element group 283: 	240 
    -- CP-element group 283: 	228 
    -- CP-element group 283: marked-predecessors 
    -- CP-element group 283: 	285 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_Sample/$entry
      -- 
    req_7439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(283), ack => WPIPE_xxconvolvexxconv_k3_2946_inst_req_0); -- 
    convolve_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(282) & convolve_CP_6526_elements(252) & convolve_CP_6526_elements(240) & convolve_CP_6526_elements(228) & convolve_CP_6526_elements(285);
      gj_convolve_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	280 
    -- CP-element group 284: 	226 
    -- CP-element group 284: 	250 
    -- CP-element group 284: 	238 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_update_start_
      -- CP-element group 284: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_Update/req
      -- CP-element group 284: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_Sample/$exit
      -- 
    ack_7440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_2946_inst_ack_0, ack => convolve_CP_6526_elements(284)); -- 
    req_7444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(284), ack => WPIPE_xxconvolvexxconv_k3_2946_inst_req_1); -- 
    -- CP-element group 285:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	317 
    -- CP-element group 285: marked-successors 
    -- CP-element group 285: 	283 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_Update/ack
      -- CP-element group 285: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_xxconvolvexxconv_k3_2946_Update/$exit
      -- 
    ack_7445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_2946_inst_ack_1, ack => convolve_CP_6526_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	108 
    -- CP-element group 286: 	127 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	288 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_Sample/req
      -- 
    req_7453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(286), ack => W_num_done_2880_delayed_1_0_2987_inst_req_0); -- 
    convolve_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(127) & convolve_CP_6526_elements(288);
      gj_convolve_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	26 
    -- CP-element group 287: marked-predecessors 
    -- CP-element group 287: 	289 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	289 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_Update/req
      -- CP-element group 287: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_update_start_
      -- 
    req_7458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(287), ack => W_num_done_2880_delayed_1_0_2987_inst_req_1); -- 
    convolve_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(289);
      gj_convolve_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: 	106 
    -- CP-element group 288: 	123 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_Sample/ack
      -- CP-element group 288: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_Sample/$exit
      -- 
    ack_7454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2880_delayed_1_0_2987_inst_ack_0, ack => convolve_CP_6526_elements(288)); -- 
    -- CP-element group 289:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	317 
    -- CP-element group 289: marked-successors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: 	29 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_Update/ack
      -- CP-element group 289: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2989_update_completed_
      -- 
    ack_7459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2880_delayed_1_0_2987_inst_ack_1, ack => convolve_CP_6526_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	108 
    -- CP-element group 290: 	127 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_sample_start_
      -- 
    req_7467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(290), ack => W_num_done_2886_delayed_1_0_2996_inst_req_0); -- 
    convolve_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(127) & convolve_CP_6526_elements(292);
      gj_convolve_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	26 
    -- CP-element group 291: marked-predecessors 
    -- CP-element group 291: 	293 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_update_start_
      -- CP-element group 291: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_Update/req
      -- 
    req_7472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(291), ack => W_num_done_2886_delayed_1_0_2996_inst_req_1); -- 
    convolve_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(26) & convolve_CP_6526_elements(293);
      gj_convolve_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	106 
    -- CP-element group 292: 	290 
    -- CP-element group 292: 	123 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_sample_completed_
      -- CP-element group 292: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_Sample/ack
      -- 
    ack_7468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2886_delayed_1_0_2996_inst_ack_0, ack => convolve_CP_6526_elements(292)); -- 
    -- CP-element group 293:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	317 
    -- CP-element group 293: marked-successors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: 	48 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_2998_Update/ack
      -- 
    ack_7473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2886_delayed_1_0_2996_inst_ack_1, ack => convolve_CP_6526_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	108 
    -- CP-element group 294: 	127 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_sample_start_
      -- CP-element group 294: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_Sample/req
      -- 
    req_7481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(294), ack => W_num_done_2891_delayed_1_0_3005_inst_req_0); -- 
    convolve_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(127) & convolve_CP_6526_elements(296);
      gj_convolve_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: marked-predecessors 
    -- CP-element group 295: 	297 
    -- CP-element group 295: 	300 
    -- CP-element group 295: 	303 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	297 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_update_start_
      -- CP-element group 295: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_Update/req
      -- 
    req_7486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(295), ack => W_num_done_2891_delayed_1_0_3005_inst_req_1); -- 
    convolve_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(297) & convolve_CP_6526_elements(300) & convolve_CP_6526_elements(303);
      gj_convolve_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	106 
    -- CP-element group 296: 	294 
    -- CP-element group 296: 	123 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_sample_completed_
      -- CP-element group 296: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_Sample/ack
      -- 
    ack_7482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2891_delayed_1_0_3005_inst_ack_0, ack => convolve_CP_6526_elements(296)); -- 
    -- CP-element group 297:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	295 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297: 	302 
    -- CP-element group 297: marked-successors 
    -- CP-element group 297: 	295 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_update_completed_
      -- CP-element group 297: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3007_Update/ack
      -- 
    ack_7487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2891_delayed_1_0_3005_inst_ack_1, ack => convolve_CP_6526_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	224 
    -- CP-element group 298: 	220 
    -- CP-element group 298: 	244 
    -- CP-element group 298: 	248 
    -- CP-element group 298: 	252 
    -- CP-element group 298: 	236 
    -- CP-element group 298: 	240 
    -- CP-element group 298: 	228 
    -- CP-element group 298: 	232 
    -- CP-element group 298: 	256 
    -- CP-element group 298: 	176 
    -- CP-element group 298: 	168 
    -- CP-element group 298: 	297 
    -- CP-element group 298: 	148 
    -- CP-element group 298: 	152 
    -- CP-element group 298: 	160 
    -- CP-element group 298: 	164 
    -- CP-element group 298: 	144 
    -- CP-element group 298: 	180 
    -- CP-element group 298: 	184 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_Sample/rr
      -- 
    rr_7495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(298), ack => type_cast_3011_inst_req_0); -- 
    convolve_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(224) & convolve_CP_6526_elements(220) & convolve_CP_6526_elements(244) & convolve_CP_6526_elements(248) & convolve_CP_6526_elements(252) & convolve_CP_6526_elements(236) & convolve_CP_6526_elements(240) & convolve_CP_6526_elements(228) & convolve_CP_6526_elements(232) & convolve_CP_6526_elements(256) & convolve_CP_6526_elements(176) & convolve_CP_6526_elements(168) & convolve_CP_6526_elements(297) & convolve_CP_6526_elements(148) & convolve_CP_6526_elements(152) & convolve_CP_6526_elements(160) & convolve_CP_6526_elements(164) & convolve_CP_6526_elements(144) & convolve_CP_6526_elements(180) & convolve_CP_6526_elements(184) & convolve_CP_6526_elements(300);
      gj_convolve_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: marked-predecessors 
    -- CP-element group 299: 	301 
    -- CP-element group 299: 	303 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	301 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_update_start_
      -- CP-element group 299: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_Update/cr
      -- 
    cr_7500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(299), ack => type_cast_3011_inst_req_1); -- 
    convolve_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(301) & convolve_CP_6526_elements(303);
      gj_convolve_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	222 
    -- CP-element group 300: 	226 
    -- CP-element group 300: 	218 
    -- CP-element group 300: 	242 
    -- CP-element group 300: 	246 
    -- CP-element group 300: 	250 
    -- CP-element group 300: 	254 
    -- CP-element group 300: 	238 
    -- CP-element group 300: 	230 
    -- CP-element group 300: 	234 
    -- CP-element group 300: 	295 
    -- CP-element group 300: 	174 
    -- CP-element group 300: 	178 
    -- CP-element group 300: 	166 
    -- CP-element group 300: 	298 
    -- CP-element group 300: 	146 
    -- CP-element group 300: 	150 
    -- CP-element group 300: 	158 
    -- CP-element group 300: 	162 
    -- CP-element group 300: 	142 
    -- CP-element group 300: 	182 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_Sample/ra
      -- 
    ra_7496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3011_inst_ack_0, ack => convolve_CP_6526_elements(300)); -- 
    -- CP-element group 301:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	299 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301: marked-successors 
    -- CP-element group 301: 	299 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3011_Update/ca
      -- 
    ca_7501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3011_inst_ack_1, ack => convolve_CP_6526_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	297 
    -- CP-element group 302: 	301 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	315 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_Sample/req
      -- 
    req_7509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(302), ack => WPIPE_output_pipe_3009_inst_req_0); -- 
    convolve_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(297) & convolve_CP_6526_elements(301) & convolve_CP_6526_elements(315) & convolve_CP_6526_elements(304);
      gj_convolve_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	295 
    -- CP-element group 303: 	299 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_update_start_
      -- CP-element group 303: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_Update/req
      -- 
    ack_7510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3009_inst_ack_0, ack => convolve_CP_6526_elements(303)); -- 
    req_7514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(303), ack => WPIPE_output_pipe_3009_inst_req_1); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	313 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3009_Update/ack
      -- 
    ack_7515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3009_inst_ack_1, ack => convolve_CP_6526_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	108 
    -- CP-element group 305: 	127 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_Sample/req
      -- 
    req_7523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(305), ack => W_num_done_2896_delayed_1_0_3013_inst_req_0); -- 
    convolve_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(108) & convolve_CP_6526_elements(127) & convolve_CP_6526_elements(307);
      gj_convolve_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	311 
    -- CP-element group 306: 	314 
    -- CP-element group 306: 	308 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_update_start_
      -- CP-element group 306: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_Update/req
      -- 
    req_7528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(306), ack => W_num_done_2896_delayed_1_0_3013_inst_req_1); -- 
    convolve_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(311) & convolve_CP_6526_elements(314) & convolve_CP_6526_elements(308);
      gj_convolve_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	106 
    -- CP-element group 307: 	123 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_Sample/ack
      -- 
    ack_7524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2896_delayed_1_0_3013_inst_ack_0, ack => convolve_CP_6526_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	313 
    -- CP-element group 308: 	309 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/assign_stmt_3015_Update/ack
      -- 
    ack_7529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2896_delayed_1_0_3013_inst_ack_1, ack => convolve_CP_6526_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	224 
    -- CP-element group 309: 	220 
    -- CP-element group 309: 	244 
    -- CP-element group 309: 	248 
    -- CP-element group 309: 	252 
    -- CP-element group 309: 	236 
    -- CP-element group 309: 	240 
    -- CP-element group 309: 	228 
    -- CP-element group 309: 	232 
    -- CP-element group 309: 	260 
    -- CP-element group 309: 	172 
    -- CP-element group 309: 	168 
    -- CP-element group 309: 	308 
    -- CP-element group 309: 	148 
    -- CP-element group 309: 	152 
    -- CP-element group 309: 	156 
    -- CP-element group 309: 	164 
    -- CP-element group 309: 	180 
    -- CP-element group 309: 	184 
    -- CP-element group 309: 	188 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_Sample/rr
      -- 
    rr_7537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(309), ack => type_cast_3019_inst_req_0); -- 
    convolve_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(224) & convolve_CP_6526_elements(220) & convolve_CP_6526_elements(244) & convolve_CP_6526_elements(248) & convolve_CP_6526_elements(252) & convolve_CP_6526_elements(236) & convolve_CP_6526_elements(240) & convolve_CP_6526_elements(228) & convolve_CP_6526_elements(232) & convolve_CP_6526_elements(260) & convolve_CP_6526_elements(172) & convolve_CP_6526_elements(168) & convolve_CP_6526_elements(308) & convolve_CP_6526_elements(148) & convolve_CP_6526_elements(152) & convolve_CP_6526_elements(156) & convolve_CP_6526_elements(164) & convolve_CP_6526_elements(180) & convolve_CP_6526_elements(184) & convolve_CP_6526_elements(188) & convolve_CP_6526_elements(311);
      gj_convolve_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	314 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_update_start_
      -- CP-element group 310: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_Update/cr
      -- 
    cr_7542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(310), ack => type_cast_3019_inst_req_1); -- 
    convolve_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(312) & convolve_CP_6526_elements(314);
      gj_convolve_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	222 
    -- CP-element group 311: 	226 
    -- CP-element group 311: 	218 
    -- CP-element group 311: 	242 
    -- CP-element group 311: 	246 
    -- CP-element group 311: 	250 
    -- CP-element group 311: 	238 
    -- CP-element group 311: 	230 
    -- CP-element group 311: 	234 
    -- CP-element group 311: 	258 
    -- CP-element group 311: 	178 
    -- CP-element group 311: 	166 
    -- CP-element group 311: 	170 
    -- CP-element group 311: 	306 
    -- CP-element group 311: 	309 
    -- CP-element group 311: 	146 
    -- CP-element group 311: 	150 
    -- CP-element group 311: 	154 
    -- CP-element group 311: 	162 
    -- CP-element group 311: 	182 
    -- CP-element group 311: 	186 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_Sample/ra
      -- 
    ra_7538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3019_inst_ack_0, ack => convolve_CP_6526_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/type_cast_3019_Update/ca
      -- 
    ca_7543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3019_inst_ack_1, ack => convolve_CP_6526_elements(312)); -- 
    -- CP-element group 313:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: 	304 
    -- CP-element group 313: 	308 
    -- CP-element group 313: marked-predecessors 
    -- CP-element group 313: 	315 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_Sample/req
      -- 
    req_7551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(313), ack => WPIPE_output_pipe_3017_inst_req_0); -- 
    convolve_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(312) & convolve_CP_6526_elements(304) & convolve_CP_6526_elements(308) & convolve_CP_6526_elements(315);
      gj_convolve_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	310 
    -- CP-element group 314: 	306 
    -- CP-element group 314:  members (6) 
      -- CP-element group 314: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_sample_completed_
      -- CP-element group 314: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_update_start_
      -- CP-element group 314: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_Sample/ack
      -- CP-element group 314: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_Update/$entry
      -- CP-element group 314: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_Update/req
      -- 
    ack_7552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3017_inst_ack_0, ack => convolve_CP_6526_elements(314)); -- 
    req_7556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(314), ack => WPIPE_output_pipe_3017_inst_req_1); -- 
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: 	302 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_update_completed_
      -- CP-element group 315: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_Update/$exit
      -- CP-element group 315: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/WPIPE_output_pipe_3017_Update/ack
      -- 
    ack_7557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3017_inst_ack_1, ack => convolve_CP_6526_elements(315)); -- 
    -- CP-element group 316:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	23 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	24 
    -- CP-element group 316:  members (1) 
      -- CP-element group 316: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_6526_elements(316) is a control-delay.
    cp_element_316_delay: control_delay_element  generic map(name => " 316_delay", delay_value => 1)  port map(req => convolve_CP_6526_elements(23), ack => convolve_CP_6526_elements(316), clk => clk, reset =>reset);
    -- CP-element group 317:  join  transition  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	285 
    -- CP-element group 317: 	271 
    -- CP-element group 317: 	278 
    -- CP-element group 317: 	216 
    -- CP-element group 317: 	289 
    -- CP-element group 317: 	293 
    -- CP-element group 317: 	26 
    -- CP-element group 317: 	315 
    -- CP-element group 317: 	209 
    -- CP-element group 317: 	202 
    -- CP-element group 317: 	195 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	20 
    -- CP-element group 317:  members (1) 
      -- CP-element group 317: 	 branch_block_stmt_2571/do_while_stmt_2588/do_while_stmt_2588_loop_body/$exit
      -- 
    convolve_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolve_CP_6526_elements(285) & convolve_CP_6526_elements(271) & convolve_CP_6526_elements(278) & convolve_CP_6526_elements(216) & convolve_CP_6526_elements(289) & convolve_CP_6526_elements(293) & convolve_CP_6526_elements(26) & convolve_CP_6526_elements(315) & convolve_CP_6526_elements(209) & convolve_CP_6526_elements(202) & convolve_CP_6526_elements(195);
      gj_convolve_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_6526_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	19 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_2571/do_while_stmt_2588/loop_exit/$exit
      -- CP-element group 318: 	 branch_block_stmt_2571/do_while_stmt_2588/loop_exit/ack
      -- 
    ack_7562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2588_branch_ack_0, ack => convolve_CP_6526_elements(318)); -- 
    -- CP-element group 319:  transition  input  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	19 
    -- CP-element group 319: successors 
    -- CP-element group 319:  members (2) 
      -- CP-element group 319: 	 branch_block_stmt_2571/do_while_stmt_2588/loop_taken/$exit
      -- CP-element group 319: 	 branch_block_stmt_2571/do_while_stmt_2588/loop_taken/ack
      -- 
    ack_7566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2588_branch_ack_1, ack => convolve_CP_6526_elements(319)); -- 
    -- CP-element group 320:  transition  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	17 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	2 
    -- CP-element group 320:  members (1) 
      -- CP-element group 320: 	 branch_block_stmt_2571/do_while_stmt_2588/$exit
      -- 
    convolve_CP_6526_elements(320) <= convolve_CP_6526_elements(17);
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	2 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_sample_completed_
      -- CP-element group 321: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_update_start_
      -- CP-element group 321: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_Sample/$exit
      -- CP-element group 321: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_Sample/ack
      -- CP-element group 321: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_Update/req
      -- 
    ack_7579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3024_inst_ack_0, ack => convolve_CP_6526_elements(321)); -- 
    req_7583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(321), ack => WPIPE_input_done_pipe_3024_inst_req_1); -- 
    -- CP-element group 322:  transition  place  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (8) 
      -- CP-element group 322: 	 branch_block_stmt_2571/assign_stmt_3026__exit__
      -- CP-element group 322: 	 branch_block_stmt_2571/loopback
      -- CP-element group 322: 	 branch_block_stmt_2571/assign_stmt_3026/$exit
      -- CP-element group 322: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_update_completed_
      -- CP-element group 322: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_Update/$exit
      -- CP-element group 322: 	 branch_block_stmt_2571/assign_stmt_3026/WPIPE_input_done_pipe_3024_Update/ack
      -- CP-element group 322: 	 branch_block_stmt_2571/loopback_PhiReq/$entry
      -- CP-element group 322: 	 branch_block_stmt_2571/loopback_PhiReq/$exit
      -- 
    ack_7584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3024_inst_ack_1, ack => convolve_CP_6526_elements(322)); -- 
    -- CP-element group 323:  merge  fork  transition  place  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: 	0 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	3 
    -- CP-element group 323: 	6 
    -- CP-element group 323: 	10 
    -- CP-element group 323: 	11 
    -- CP-element group 323: 	14 
    -- CP-element group 323:  members (22) 
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_update_start_
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_Update/cr
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_Sample/rr
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2586_Update/cr
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_size_pipe_2584_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_2571/merge_stmt_2572__exit__
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587__entry__
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/$entry
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_update_start_
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/RPIPE_num_out_pipe_2574_Sample/rr
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2576_Update/cr
      -- CP-element group 323: 	 branch_block_stmt_2571/assign_stmt_2577_to_assign_stmt_2587/SUB_u16_u16_2581_update_start_
      -- CP-element group 323: 	 branch_block_stmt_2571/merge_stmt_2572_PhiReqMerge
      -- CP-element group 323: 	 branch_block_stmt_2571/merge_stmt_2572_PhiAck/$entry
      -- CP-element group 323: 	 branch_block_stmt_2571/merge_stmt_2572_PhiAck/$exit
      -- CP-element group 323: 	 branch_block_stmt_2571/merge_stmt_2572_PhiAck/dummy
      -- 
    cr_6600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(323), ack => SUB_u16_u16_2581_inst_req_1); -- 
    rr_6613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(323), ack => RPIPE_size_pipe_2584_inst_req_0); -- 
    cr_6628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(323), ack => SUB_u16_u16_2586_inst_req_1); -- 
    rr_6557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(323), ack => RPIPE_num_out_pipe_2574_inst_req_0); -- 
    cr_6572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_6526_elements(323), ack => SUB_u16_u16_2576_inst_req_1); -- 
    convolve_CP_6526_elements(323) <= OrReduce(convolve_CP_6526_elements(322) & convolve_CP_6526_elements(0));
    convolve_do_while_stmt_2588_terminator_7567: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_2588_terminator_7567", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_6526_elements(20),loop_continue => convolve_CP_6526_elements(319),loop_terminate => convolve_CP_6526_elements(318),loop_back => convolve_CP_6526_elements(18),loop_exit => convolve_CP_6526_elements(17),clk => clk, reset => reset); -- 
    phi_stmt_2590_phi_seq_6693_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6526_elements(37);
      convolve_CP_6526_elements(40)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6526_elements(40);
      convolve_CP_6526_elements(41)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6526_elements(42);
      convolve_CP_6526_elements(38) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6526_elements(35);
      convolve_CP_6526_elements(44)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6526_elements(46);
      convolve_CP_6526_elements(45)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6526_elements(47);
      convolve_CP_6526_elements(36) <= phi_mux_reqs(1);
      phi_stmt_2590_phi_seq_6693 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2590_phi_seq_6693") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6526_elements(31), 
          phi_sample_ack => convolve_CP_6526_elements(32), 
          phi_update_req => convolve_CP_6526_elements(33), 
          phi_update_ack => convolve_CP_6526_elements(34), 
          phi_mux_ack => convolve_CP_6526_elements(39), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2596_phi_seq_6737_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6526_elements(56);
      convolve_CP_6526_elements(59)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6526_elements(59);
      convolve_CP_6526_elements(60)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6526_elements(61);
      convolve_CP_6526_elements(57) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6526_elements(54);
      convolve_CP_6526_elements(63)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6526_elements(65);
      convolve_CP_6526_elements(64)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6526_elements(66);
      convolve_CP_6526_elements(55) <= phi_mux_reqs(1);
      phi_stmt_2596_phi_seq_6737 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2596_phi_seq_6737") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6526_elements(50), 
          phi_sample_ack => convolve_CP_6526_elements(51), 
          phi_update_req => convolve_CP_6526_elements(52), 
          phi_update_ack => convolve_CP_6526_elements(53), 
          phi_mux_ack => convolve_CP_6526_elements(58), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2601_phi_seq_6781_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6526_elements(75);
      convolve_CP_6526_elements(78)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6526_elements(78);
      convolve_CP_6526_elements(79)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6526_elements(80);
      convolve_CP_6526_elements(76) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6526_elements(73);
      convolve_CP_6526_elements(82)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6526_elements(84);
      convolve_CP_6526_elements(83)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6526_elements(85);
      convolve_CP_6526_elements(74) <= phi_mux_reqs(1);
      phi_stmt_2601_phi_seq_6781 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2601_phi_seq_6781") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6526_elements(69), 
          phi_sample_ack => convolve_CP_6526_elements(70), 
          phi_update_req => convolve_CP_6526_elements(71), 
          phi_update_ack => convolve_CP_6526_elements(72), 
          phi_mux_ack => convolve_CP_6526_elements(77), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2606_phi_seq_6825_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6526_elements(94);
      convolve_CP_6526_elements(97)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6526_elements(97);
      convolve_CP_6526_elements(98)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6526_elements(99);
      convolve_CP_6526_elements(95) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6526_elements(92);
      convolve_CP_6526_elements(101)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6526_elements(103);
      convolve_CP_6526_elements(102)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6526_elements(104);
      convolve_CP_6526_elements(93) <= phi_mux_reqs(1);
      phi_stmt_2606_phi_seq_6825 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2606_phi_seq_6825") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6526_elements(88), 
          phi_sample_ack => convolve_CP_6526_elements(89), 
          phi_update_req => convolve_CP_6526_elements(90), 
          phi_update_ack => convolve_CP_6526_elements(91), 
          phi_mux_ack => convolve_CP_6526_elements(96), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2611_phi_seq_6869_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6526_elements(111);
      convolve_CP_6526_elements(114)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6526_elements(114);
      convolve_CP_6526_elements(115)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6526_elements(116);
      convolve_CP_6526_elements(112) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6526_elements(109);
      convolve_CP_6526_elements(118)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6526_elements(120);
      convolve_CP_6526_elements(119)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6526_elements(121);
      convolve_CP_6526_elements(110) <= phi_mux_reqs(1);
      phi_stmt_2611_phi_seq_6869 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2611_phi_seq_6869") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6526_elements(25), 
          phi_sample_ack => convolve_CP_6526_elements(107), 
          phi_update_req => convolve_CP_6526_elements(27), 
          phi_update_ack => convolve_CP_6526_elements(108), 
          phi_mux_ack => convolve_CP_6526_elements(113), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2617_phi_seq_6913_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_6526_elements(130);
      convolve_CP_6526_elements(133)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_6526_elements(133);
      convolve_CP_6526_elements(134)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_6526_elements(135);
      convolve_CP_6526_elements(131) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_6526_elements(128);
      convolve_CP_6526_elements(137)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_6526_elements(139);
      convolve_CP_6526_elements(138)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_6526_elements(140);
      convolve_CP_6526_elements(129) <= phi_mux_reqs(1);
      phi_stmt_2617_phi_seq_6913 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2617_phi_seq_6913") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_6526_elements(124), 
          phi_sample_ack => convolve_CP_6526_elements(125), 
          phi_update_req => convolve_CP_6526_elements(126), 
          phi_update_ack => convolve_CP_6526_elements(127), 
          phi_mux_ack => convolve_CP_6526_elements(132), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6645_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_6526_elements(21);
        preds(1)  <= convolve_CP_6526_elements(22);
        entry_tmerge_6645 : transition_merge -- 
          generic map(name => " entry_tmerge_6645")
          port map (preds => preds, symbol_out => convolve_CP_6526_elements(23));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_i16_i16_2867_wire : std_logic_vector(15 downto 0);
    signal ADD_i16_i16_2870_wire : std_logic_vector(15 downto 0);
    signal ADD_i16_i16_2879_wire : std_logic_vector(15 downto 0);
    signal ADD_i16_i16_2882_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2954_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2974_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2983_wire : std_logic_vector(15 downto 0);
    signal ADD_u2_u2_2963_wire : std_logic_vector(1 downto 0);
    signal AND_u1_u1_2920_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2626_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2756_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2759_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2629_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2893_wire : std_logic_vector(0 downto 0);
    signal MUL_i16_i16_2828_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2834_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2840_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2846_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2852_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2858_wire : std_logic_vector(15 downto 0);
    signal MUX_2964_wire : std_logic_vector(1 downto 0);
    signal MUX_2975_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_3023_wire : std_logic_vector(0 downto 0);
    signal RPIPE_num_out_pipe_2574_wire : std_logic_vector(15 downto 0);
    signal RPIPE_num_out_pipe_2579_wire : std_logic_vector(15 downto 0);
    signal RPIPE_size_pipe_2584_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_2815_2815_delayed_1_0_2911 : std_logic_vector(15 downto 0);
    signal UGT_u2_u1_2706_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_2703_wire : std_logic_vector(0 downto 0);
    signal acc1_2590 : std_logic_vector(15 downto 0);
    signal acc1_2772_delayed_1_0_2863 : std_logic_vector(15 downto 0);
    signal acc2_2596 : std_logic_vector(15 downto 0);
    signal acc2_2781_delayed_1_0_2875 : std_logic_vector(15 downto 0);
    signal acc_val1_2872 : std_logic_vector(15 downto 0);
    signal acc_val2_2884 : std_logic_vector(15 downto 0);
    signal all_done_flag_2927 : std_logic_vector(0 downto 0);
    signal chl_2617 : std_logic_vector(15 downto 0);
    signal chl_done_2889 : std_logic_vector(0 downto 0);
    signal col_2606 : std_logic_vector(15 downto 0);
    signal col_done_2901 : std_logic_vector(0 downto 0);
    signal iread1_2672 : std_logic_vector(15 downto 0);
    signal iread2_2681 : std_logic_vector(15 downto 0);
    signal iread3_2690 : std_logic_vector(15 downto 0);
    signal iread4_2699 : std_logic_vector(15 downto 0);
    signal ival1_2740 : std_logic_vector(15 downto 0);
    signal ival2_2744 : std_logic_vector(15 downto 0);
    signal ival3_2748 : std_logic_vector(15 downto 0);
    signal ival4_2752 : std_logic_vector(15 downto 0);
    signal konst_2575_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2580_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2585_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2625_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2628_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2705_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2755_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2758_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2892_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2909_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2951_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2953_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2960_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2962_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2971_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2973_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2982_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2992_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3001_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3025_wire_constant : std_logic_vector(7 downto 0);
    signal kread1_2794 : std_logic_vector(15 downto 0);
    signal kread2_2803 : std_logic_vector(15 downto 0);
    signal kread3_2812 : std_logic_vector(15 downto 0);
    signal kval1_2816 : std_logic_vector(15 downto 0);
    signal kval2_2820 : std_logic_vector(15 downto 0);
    signal kval3_2824 : std_logic_vector(15 downto 0);
    signal mul_val1_2830 : std_logic_vector(15 downto 0);
    signal mul_val2_2836 : std_logic_vector(15 downto 0);
    signal mul_val3_2842 : std_logic_vector(15 downto 0);
    signal mul_val4_2848 : std_logic_vector(15 downto 0);
    signal mul_val5_2854 : std_logic_vector(15 downto 0);
    signal mul_val6_2860 : std_logic_vector(15 downto 0);
    signal n_chl_2956 : std_logic_vector(15 downto 0);
    signal n_chl_2956_2621_buffered : std_logic_vector(15 downto 0);
    signal n_col_2978 : std_logic_vector(15 downto 0);
    signal n_col_2978_2610_buffered : std_logic_vector(15 downto 0);
    signal n_num_2967 : std_logic_vector(1 downto 0);
    signal n_num_2967_2616_buffered : std_logic_vector(1 downto 0);
    signal n_row_2986 : std_logic_vector(15 downto 0);
    signal n_row_2986_2605_buffered : std_logic_vector(15 downto 0);
    signal nacc1_2995 : std_logic_vector(15 downto 0);
    signal nacc1_2995_2595_buffered : std_logic_vector(15 downto 0);
    signal nacc2_3004 : std_logic_vector(15 downto 0);
    signal nacc2_3004_2600_buffered : std_logic_vector(15 downto 0);
    signal num_2611 : std_logic_vector(1 downto 0);
    signal num_chl_2587 : std_logic_vector(15 downto 0);
    signal num_col_2582 : std_logic_vector(15 downto 0);
    signal num_done_2880_delayed_1_0_2989 : std_logic_vector(0 downto 0);
    signal num_done_2886_delayed_1_0_2998 : std_logic_vector(0 downto 0);
    signal num_done_2891_delayed_1_0_3007 : std_logic_vector(0 downto 0);
    signal num_done_2896 : std_logic_vector(0 downto 0);
    signal num_done_2896_delayed_1_0_3015 : std_logic_vector(0 downto 0);
    signal num_row_2577 : std_logic_vector(15 downto 0);
    signal out_done_flag_2916 : std_logic_vector(0 downto 0);
    signal read_ip_2608_delayed_1_0_2666 : std_logic_vector(0 downto 0);
    signal read_ip_2614_delayed_1_0_2675 : std_logic_vector(0 downto 0);
    signal read_ip_2620_delayed_1_0_2684 : std_logic_vector(0 downto 0);
    signal read_ip_2626_delayed_1_0_2693 : std_logic_vector(0 downto 0);
    signal read_ip_2631 : std_logic_vector(0 downto 0);
    signal read_k_2706_delayed_1_0_2788 : std_logic_vector(0 downto 0);
    signal read_k_2712_delayed_1_0_2797 : std_logic_vector(0 downto 0);
    signal read_k_2718_delayed_1_0_2806 : std_logic_vector(0 downto 0);
    signal read_k_2761 : std_logic_vector(0 downto 0);
    signal row_2601 : std_logic_vector(15 downto 0);
    signal row_done_2906 : std_logic_vector(0 downto 0);
    signal store_kernel_2829_delayed_1_0_2930 : std_logic_vector(0 downto 0);
    signal store_kernel_2833_delayed_1_0_2937 : std_logic_vector(0 downto 0);
    signal store_kernel_2837_delayed_1_0_2944 : std_logic_vector(0 downto 0);
    signal store_kernel_2922 : std_logic_vector(0 downto 0);
    signal temp1_1_2651 : std_logic_vector(15 downto 0);
    signal temp1_2_2655 : std_logic_vector(15 downto 0);
    signal temp1_3_2659 : std_logic_vector(15 downto 0);
    signal temp1_4_2663 : std_logic_vector(15 downto 0);
    signal temp2_1_2635 : std_logic_vector(15 downto 0);
    signal temp2_2_2639 : std_logic_vector(15 downto 0);
    signal temp2_3_2643 : std_logic_vector(15 downto 0);
    signal temp2_4_2647 : std_logic_vector(15 downto 0);
    signal tempk1_1_2765 : std_logic_vector(15 downto 0);
    signal tempk1_2_2769 : std_logic_vector(15 downto 0);
    signal tempk1_3_2773 : std_logic_vector(15 downto 0);
    signal tempk2_1_2777 : std_logic_vector(15 downto 0);
    signal tempk2_2_2781 : std_logic_vector(15 downto 0);
    signal tempk2_3_2785 : std_logic_vector(15 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2599_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2604_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2609_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2615_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_2620_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3011_wire : std_logic_vector(15 downto 0);
    signal type_cast_3019_wire : std_logic_vector(15 downto 0);
    signal write_input_2640_delayed_1_0_2711 : std_logic_vector(0 downto 0);
    signal write_input_2644_delayed_1_0_2718 : std_logic_vector(0 downto 0);
    signal write_input_2648_delayed_1_0_2725 : std_logic_vector(0 downto 0);
    signal write_input_2652_delayed_1_0_2732 : std_logic_vector(0 downto 0);
    signal write_input_2708 : std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip4
    signal xxconvolvexxconv_ip4_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip4_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip4_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip4
    signal xxconvolvexxconv_ip4_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip4_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip4_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_2575_wire_constant <= "0000000000000001";
    konst_2580_wire_constant <= "0000000000000001";
    konst_2585_wire_constant <= "0000000000000001";
    konst_2625_wire_constant <= "0000000000000000";
    konst_2628_wire_constant <= "10";
    konst_2705_wire_constant <= "00";
    konst_2755_wire_constant <= "0000000000000000";
    konst_2758_wire_constant <= "0000000000000000";
    konst_2892_wire_constant <= "10";
    konst_2909_wire_constant <= "0000000000000001";
    konst_2951_wire_constant <= "0000000000000000";
    konst_2953_wire_constant <= "0000000000000001";
    konst_2960_wire_constant <= "00";
    konst_2962_wire_constant <= "01";
    konst_2971_wire_constant <= "0000000000000000";
    konst_2973_wire_constant <= "0000000000000001";
    konst_2982_wire_constant <= "0000000000000010";
    konst_2992_wire_constant <= "0000000000000000";
    konst_3001_wire_constant <= "0000000000000000";
    konst_3025_wire_constant <= "00000001";
    type_cast_2594_wire_constant <= "0000000000000000";
    type_cast_2599_wire_constant <= "0000000000000000";
    type_cast_2604_wire_constant <= "0000000000000000";
    type_cast_2609_wire_constant <= "0000000000000000";
    type_cast_2615_wire_constant <= "00";
    type_cast_2620_wire_constant <= "0000000000000000";
    phi_stmt_2590: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2594_wire_constant & nacc1_2995_2595_buffered;
      req <= phi_stmt_2590_req_0 & phi_stmt_2590_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2590",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2590_ack_0,
          idata => idata,
          odata => acc1_2590,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2590
    phi_stmt_2596: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2599_wire_constant & nacc2_3004_2600_buffered;
      req <= phi_stmt_2596_req_0 & phi_stmt_2596_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2596",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2596_ack_0,
          idata => idata,
          odata => acc2_2596,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2596
    phi_stmt_2601: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2604_wire_constant & n_row_2986_2605_buffered;
      req <= phi_stmt_2601_req_0 & phi_stmt_2601_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2601",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2601_ack_0,
          idata => idata,
          odata => row_2601,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2601
    phi_stmt_2606: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2609_wire_constant & n_col_2978_2610_buffered;
      req <= phi_stmt_2606_req_0 & phi_stmt_2606_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2606",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2606_ack_0,
          idata => idata,
          odata => col_2606,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2606
    phi_stmt_2611: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2615_wire_constant & n_num_2967_2616_buffered;
      req <= phi_stmt_2611_req_0 & phi_stmt_2611_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2611",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2611_ack_0,
          idata => idata,
          odata => num_2611,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2611
    phi_stmt_2617: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2620_wire_constant & n_chl_2956_2621_buffered;
      req <= phi_stmt_2617_req_0 & phi_stmt_2617_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2617",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2617_ack_0,
          idata => idata,
          odata => chl_2617,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2617
    -- flow-through select operator MUX_2671_inst
    iread1_2672 <= temp2_1_2635 when (read_ip_2608_delayed_1_0_2666(0) /=  '0') else temp1_1_2651;
    -- flow-through select operator MUX_2680_inst
    iread2_2681 <= temp2_2_2639 when (read_ip_2614_delayed_1_0_2675(0) /=  '0') else temp1_2_2655;
    -- flow-through select operator MUX_2689_inst
    iread3_2690 <= temp2_3_2643 when (read_ip_2620_delayed_1_0_2684(0) /=  '0') else temp1_3_2659;
    -- flow-through select operator MUX_2698_inst
    iread4_2699 <= temp2_4_2647 when (read_ip_2626_delayed_1_0_2693(0) /=  '0') else temp1_4_2663;
    -- flow-through select operator MUX_2793_inst
    kread1_2794 <= tempk1_1_2765 when (read_k_2706_delayed_1_0_2788(0) /=  '0') else tempk2_1_2777;
    -- flow-through select operator MUX_2802_inst
    kread2_2803 <= tempk1_2_2769 when (read_k_2712_delayed_1_0_2797(0) /=  '0') else tempk2_2_2781;
    -- flow-through select operator MUX_2811_inst
    kread3_2812 <= tempk1_3_2773 when (read_k_2718_delayed_1_0_2806(0) /=  '0') else tempk2_3_2785;
    -- flow-through select operator MUX_2955_inst
    n_chl_2956 <= konst_2951_wire_constant when (chl_done_2889(0) /=  '0') else ADD_u16_u16_2954_wire;
    -- flow-through select operator MUX_2964_inst
    MUX_2964_wire <= konst_2960_wire_constant when (num_done_2896(0) /=  '0') else ADD_u2_u2_2963_wire;
    -- flow-through select operator MUX_2966_inst
    n_num_2967 <= MUX_2964_wire when (chl_done_2889(0) /=  '0') else num_2611;
    -- flow-through select operator MUX_2975_inst
    MUX_2975_wire <= konst_2971_wire_constant when (col_done_2901(0) /=  '0') else ADD_u16_u16_2974_wire;
    -- flow-through select operator MUX_2977_inst
    n_col_2978 <= MUX_2975_wire when (num_done_2896(0) /=  '0') else col_2606;
    -- flow-through select operator MUX_2985_inst
    n_row_2986 <= ADD_u16_u16_2983_wire when (row_done_2906(0) /=  '0') else row_2601;
    -- flow-through select operator MUX_2994_inst
    nacc1_2995 <= konst_2992_wire_constant when (num_done_2880_delayed_1_0_2989(0) /=  '0') else acc_val1_2872;
    -- flow-through select operator MUX_3003_inst
    nacc2_3004 <= konst_3001_wire_constant when (num_done_2886_delayed_1_0_2998(0) /=  '0') else acc_val2_2884;
    W_acc1_2772_delayed_1_0_2861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc1_2772_delayed_1_0_2861_inst_req_0;
      W_acc1_2772_delayed_1_0_2861_inst_ack_0<= wack(0);
      rreq(0) <= W_acc1_2772_delayed_1_0_2861_inst_req_1;
      W_acc1_2772_delayed_1_0_2861_inst_ack_1<= rack(0);
      W_acc1_2772_delayed_1_0_2861_inst : InterlockBuffer generic map ( -- 
        name => "W_acc1_2772_delayed_1_0_2861_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc1_2590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc1_2772_delayed_1_0_2863,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_acc2_2781_delayed_1_0_2873_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc2_2781_delayed_1_0_2873_inst_req_0;
      W_acc2_2781_delayed_1_0_2873_inst_ack_0<= wack(0);
      rreq(0) <= W_acc2_2781_delayed_1_0_2873_inst_req_1;
      W_acc2_2781_delayed_1_0_2873_inst_ack_1<= rack(0);
      W_acc2_2781_delayed_1_0_2873_inst : InterlockBuffer generic map ( -- 
        name => "W_acc2_2781_delayed_1_0_2873_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc2_2596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc2_2781_delayed_1_0_2875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2880_delayed_1_0_2987_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2880_delayed_1_0_2987_inst_req_0;
      W_num_done_2880_delayed_1_0_2987_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2880_delayed_1_0_2987_inst_req_1;
      W_num_done_2880_delayed_1_0_2987_inst_ack_1<= rack(0);
      W_num_done_2880_delayed_1_0_2987_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2880_delayed_1_0_2987_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2896,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2880_delayed_1_0_2989,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2886_delayed_1_0_2996_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2886_delayed_1_0_2996_inst_req_0;
      W_num_done_2886_delayed_1_0_2996_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2886_delayed_1_0_2996_inst_req_1;
      W_num_done_2886_delayed_1_0_2996_inst_ack_1<= rack(0);
      W_num_done_2886_delayed_1_0_2996_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2886_delayed_1_0_2996_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2896,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2886_delayed_1_0_2998,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2891_delayed_1_0_3005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2891_delayed_1_0_3005_inst_req_0;
      W_num_done_2891_delayed_1_0_3005_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2891_delayed_1_0_3005_inst_req_1;
      W_num_done_2891_delayed_1_0_3005_inst_ack_1<= rack(0);
      W_num_done_2891_delayed_1_0_3005_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2891_delayed_1_0_3005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2896,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2891_delayed_1_0_3007,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2896_delayed_1_0_3013_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2896_delayed_1_0_3013_inst_req_0;
      W_num_done_2896_delayed_1_0_3013_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2896_delayed_1_0_3013_inst_req_1;
      W_num_done_2896_delayed_1_0_3013_inst_ack_1<= rack(0);
      W_num_done_2896_delayed_1_0_3013_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2896_delayed_1_0_3013_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2896,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2896_delayed_1_0_3015,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2608_delayed_1_0_2664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2608_delayed_1_0_2664_inst_req_0;
      W_read_ip_2608_delayed_1_0_2664_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2608_delayed_1_0_2664_inst_req_1;
      W_read_ip_2608_delayed_1_0_2664_inst_ack_1<= rack(0);
      W_read_ip_2608_delayed_1_0_2664_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2608_delayed_1_0_2664_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2608_delayed_1_0_2666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2614_delayed_1_0_2673_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2614_delayed_1_0_2673_inst_req_0;
      W_read_ip_2614_delayed_1_0_2673_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2614_delayed_1_0_2673_inst_req_1;
      W_read_ip_2614_delayed_1_0_2673_inst_ack_1<= rack(0);
      W_read_ip_2614_delayed_1_0_2673_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2614_delayed_1_0_2673_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2614_delayed_1_0_2675,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2620_delayed_1_0_2682_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2620_delayed_1_0_2682_inst_req_0;
      W_read_ip_2620_delayed_1_0_2682_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2620_delayed_1_0_2682_inst_req_1;
      W_read_ip_2620_delayed_1_0_2682_inst_ack_1<= rack(0);
      W_read_ip_2620_delayed_1_0_2682_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2620_delayed_1_0_2682_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2620_delayed_1_0_2684,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_2626_delayed_1_0_2691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_2626_delayed_1_0_2691_inst_req_0;
      W_read_ip_2626_delayed_1_0_2691_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_2626_delayed_1_0_2691_inst_req_1;
      W_read_ip_2626_delayed_1_0_2691_inst_ack_1<= rack(0);
      W_read_ip_2626_delayed_1_0_2691_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_2626_delayed_1_0_2691_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_2631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_2626_delayed_1_0_2693,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2706_delayed_1_0_2786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2706_delayed_1_0_2786_inst_req_0;
      W_read_k_2706_delayed_1_0_2786_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2706_delayed_1_0_2786_inst_req_1;
      W_read_k_2706_delayed_1_0_2786_inst_ack_1<= rack(0);
      W_read_k_2706_delayed_1_0_2786_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2706_delayed_1_0_2786_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2706_delayed_1_0_2788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2712_delayed_1_0_2795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2712_delayed_1_0_2795_inst_req_0;
      W_read_k_2712_delayed_1_0_2795_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2712_delayed_1_0_2795_inst_req_1;
      W_read_k_2712_delayed_1_0_2795_inst_ack_1<= rack(0);
      W_read_k_2712_delayed_1_0_2795_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2712_delayed_1_0_2795_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2712_delayed_1_0_2797,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2718_delayed_1_0_2804_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2718_delayed_1_0_2804_inst_req_0;
      W_read_k_2718_delayed_1_0_2804_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2718_delayed_1_0_2804_inst_req_1;
      W_read_k_2718_delayed_1_0_2804_inst_ack_1<= rack(0);
      W_read_k_2718_delayed_1_0_2804_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2718_delayed_1_0_2804_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2718_delayed_1_0_2806,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2829_delayed_1_0_2928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2829_delayed_1_0_2928_inst_req_0;
      W_store_kernel_2829_delayed_1_0_2928_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2829_delayed_1_0_2928_inst_req_1;
      W_store_kernel_2829_delayed_1_0_2928_inst_ack_1<= rack(0);
      W_store_kernel_2829_delayed_1_0_2928_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2829_delayed_1_0_2928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2829_delayed_1_0_2930,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2833_delayed_1_0_2935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2833_delayed_1_0_2935_inst_req_0;
      W_store_kernel_2833_delayed_1_0_2935_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2833_delayed_1_0_2935_inst_req_1;
      W_store_kernel_2833_delayed_1_0_2935_inst_ack_1<= rack(0);
      W_store_kernel_2833_delayed_1_0_2935_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2833_delayed_1_0_2935_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2833_delayed_1_0_2937,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2837_delayed_1_0_2942_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2837_delayed_1_0_2942_inst_req_0;
      W_store_kernel_2837_delayed_1_0_2942_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2837_delayed_1_0_2942_inst_req_1;
      W_store_kernel_2837_delayed_1_0_2942_inst_ack_1<= rack(0);
      W_store_kernel_2837_delayed_1_0_2942_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2837_delayed_1_0_2942_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2837_delayed_1_0_2944,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2640_delayed_1_0_2709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2640_delayed_1_0_2709_inst_req_0;
      W_write_input_2640_delayed_1_0_2709_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2640_delayed_1_0_2709_inst_req_1;
      W_write_input_2640_delayed_1_0_2709_inst_ack_1<= rack(0);
      W_write_input_2640_delayed_1_0_2709_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2640_delayed_1_0_2709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2640_delayed_1_0_2711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2644_delayed_1_0_2716_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2644_delayed_1_0_2716_inst_req_0;
      W_write_input_2644_delayed_1_0_2716_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2644_delayed_1_0_2716_inst_req_1;
      W_write_input_2644_delayed_1_0_2716_inst_ack_1<= rack(0);
      W_write_input_2644_delayed_1_0_2716_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2644_delayed_1_0_2716_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2644_delayed_1_0_2718,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2648_delayed_1_0_2723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2648_delayed_1_0_2723_inst_req_0;
      W_write_input_2648_delayed_1_0_2723_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2648_delayed_1_0_2723_inst_req_1;
      W_write_input_2648_delayed_1_0_2723_inst_ack_1<= rack(0);
      W_write_input_2648_delayed_1_0_2723_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2648_delayed_1_0_2723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2648_delayed_1_0_2725,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_2652_delayed_1_0_2730_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_2652_delayed_1_0_2730_inst_req_0;
      W_write_input_2652_delayed_1_0_2730_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_2652_delayed_1_0_2730_inst_req_1;
      W_write_input_2652_delayed_1_0_2730_inst_ack_1<= rack(0);
      W_write_input_2652_delayed_1_0_2730_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_2652_delayed_1_0_2730_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_2652_delayed_1_0_2732,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_2956_2621_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_2956_2621_buf_req_0;
      n_chl_2956_2621_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_2956_2621_buf_req_1;
      n_chl_2956_2621_buf_ack_1<= rack(0);
      n_chl_2956_2621_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_2956_2621_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_2956,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_2956_2621_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_2978_2610_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_2978_2610_buf_req_0;
      n_col_2978_2610_buf_ack_0<= wack(0);
      rreq(0) <= n_col_2978_2610_buf_req_1;
      n_col_2978_2610_buf_ack_1<= rack(0);
      n_col_2978_2610_buf : InterlockBuffer generic map ( -- 
        name => "n_col_2978_2610_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_2978,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_2978_2610_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_num_2967_2616_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_num_2967_2616_buf_req_0;
      n_num_2967_2616_buf_ack_0<= wack(0);
      rreq(0) <= n_num_2967_2616_buf_req_1;
      n_num_2967_2616_buf_ack_1<= rack(0);
      n_num_2967_2616_buf : InterlockBuffer generic map ( -- 
        name => "n_num_2967_2616_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_num_2967,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_num_2967_2616_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_2986_2605_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_2986_2605_buf_req_0;
      n_row_2986_2605_buf_ack_0<= wack(0);
      rreq(0) <= n_row_2986_2605_buf_req_1;
      n_row_2986_2605_buf_ack_1<= rack(0);
      n_row_2986_2605_buf : InterlockBuffer generic map ( -- 
        name => "n_row_2986_2605_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_2986,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_2986_2605_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc1_2995_2595_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc1_2995_2595_buf_req_0;
      nacc1_2995_2595_buf_ack_0<= wack(0);
      rreq(0) <= nacc1_2995_2595_buf_req_1;
      nacc1_2995_2595_buf_ack_1<= rack(0);
      nacc1_2995_2595_buf : InterlockBuffer generic map ( -- 
        name => "nacc1_2995_2595_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc1_2995,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc1_2995_2595_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc2_3004_2600_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc2_3004_2600_buf_req_0;
      nacc2_3004_2600_buf_ack_0<= wack(0);
      rreq(0) <= nacc2_3004_2600_buf_req_1;
      nacc2_3004_2600_buf_ack_1<= rack(0);
      nacc2_3004_2600_buf : InterlockBuffer generic map ( -- 
        name => "nacc2_3004_2600_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc2_3004,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc2_3004_2600_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2739_inst
    process(iread1_2672) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread1_2672(15 downto 0);
      ival1_2740 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2743_inst
    process(iread2_2681) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread2_2681(15 downto 0);
      ival2_2744 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2747_inst
    process(iread3_2690) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread3_2690(15 downto 0);
      ival3_2748 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2751_inst
    process(iread4_2699) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread4_2699(15 downto 0);
      ival4_2752 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2815_inst
    process(kread1_2794) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread1_2794(15 downto 0);
      kval1_2816 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2819_inst
    process(kread2_2803) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread2_2803(15 downto 0);
      kval2_2820 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2823_inst
    process(kread3_2812) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread3_2812(15 downto 0);
      kval3_2824 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2829_inst
    process(MUL_i16_i16_2828_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2828_wire(15 downto 0);
      mul_val1_2830 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2835_inst
    process(MUL_i16_i16_2834_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2834_wire(15 downto 0);
      mul_val2_2836 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2841_inst
    process(MUL_i16_i16_2840_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2840_wire(15 downto 0);
      mul_val3_2842 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2847_inst
    process(MUL_i16_i16_2846_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2846_wire(15 downto 0);
      mul_val4_2848 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2853_inst
    process(MUL_i16_i16_2852_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2852_wire(15 downto 0);
      mul_val5_2854 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2859_inst
    process(MUL_i16_i16_2858_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2858_wire(15 downto 0);
      mul_val6_2860 <= tmp_var; -- 
    end process;
    type_cast_3011_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_3011_inst_req_0;
      type_cast_3011_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_3011_inst_req_1;
      type_cast_3011_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  num_done_2891_delayed_1_0_3007(0);
      type_cast_3011_inst_gI: SplitGuardInterface generic map(name => "type_cast_3011_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_3011_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3011_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val1_2872,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3011_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_3019_inst_req_0;
      type_cast_3019_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_3019_inst_req_1;
      type_cast_3019_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  num_done_2896_delayed_1_0_3015(0);
      type_cast_3019_inst_gI: SplitGuardInterface generic map(name => "type_cast_3019_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_3019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val2_2884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3019_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_2588_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_3023_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2588_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2588_branch_req_0,
          ack0 => do_while_stmt_2588_branch_ack_0,
          ack1 => do_while_stmt_2588_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_2867_inst
    process(acc1_2772_delayed_1_0_2863, mul_val1_2830) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc1_2772_delayed_1_0_2863, mul_val1_2830, tmp_var);
      ADD_i16_i16_2867_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2870_inst
    process(mul_val2_2836, mul_val3_2842) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val2_2836, mul_val3_2842, tmp_var);
      ADD_i16_i16_2870_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2871_inst
    process(ADD_i16_i16_2867_wire, ADD_i16_i16_2870_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i16_i16_2867_wire, ADD_i16_i16_2870_wire, tmp_var);
      acc_val1_2872 <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2879_inst
    process(acc2_2781_delayed_1_0_2875, mul_val4_2848) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc2_2781_delayed_1_0_2875, mul_val4_2848, tmp_var);
      ADD_i16_i16_2879_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2882_inst
    process(mul_val5_2854, mul_val6_2860) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_2854, mul_val6_2860, tmp_var);
      ADD_i16_i16_2882_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2883_inst
    process(ADD_i16_i16_2879_wire, ADD_i16_i16_2882_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i16_i16_2879_wire, ADD_i16_i16_2882_wire, tmp_var);
      acc_val2_2884 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2954_inst
    process(chl_2617) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_2617, konst_2953_wire_constant, tmp_var);
      ADD_u16_u16_2954_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2974_inst
    process(col_2606) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_2606, konst_2973_wire_constant, tmp_var);
      ADD_u16_u16_2974_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2983_inst
    process(row_2601) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_2601, konst_2982_wire_constant, tmp_var);
      ADD_u16_u16_2983_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u2_u2_2963_inst
    process(num_2611) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_2611, konst_2962_wire_constant, tmp_var);
      ADD_u2_u2_2963_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2707_inst
    process(ULT_u16_u1_2703_wire, UGT_u2_u1_2706_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ULT_u16_u1_2703_wire, UGT_u2_u1_2706_wire, tmp_var);
      write_input_2708 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2760_inst
    process(EQ_u16_u1_2756_wire, EQ_u16_u1_2759_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u16_u1_2756_wire, EQ_u16_u1_2759_wire, tmp_var);
      read_k_2761 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2895_inst
    process(EQ_u2_u1_2893_wire, chl_done_2889) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_2893_wire, chl_done_2889, tmp_var);
      num_done_2896 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2905_inst
    process(col_done_2901, num_done_2896) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_2901, num_done_2896, tmp_var);
      row_done_2906 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2920_inst
    process(out_done_flag_2916, col_done_2901) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2916, col_done_2901, tmp_var);
      AND_u1_u1_2920_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2926_inst
    process(out_done_flag_2916, row_done_2906) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2916, row_done_2906, tmp_var);
      all_done_flag_2927 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2626_inst
    process(col_2606) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2606, konst_2625_wire_constant, tmp_var);
      EQ_u16_u1_2626_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2756_inst
    process(col_2606) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2606, konst_2755_wire_constant, tmp_var);
      EQ_u16_u1_2756_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2759_inst
    process(row_2601) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(row_2601, konst_2758_wire_constant, tmp_var);
      EQ_u16_u1_2759_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2888_inst
    process(chl_2617, num_chl_2587) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(chl_2617, num_chl_2587, tmp_var);
      chl_done_2889 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2900_inst
    process(col_2606, num_col_2582) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_2606, num_col_2582, tmp_var);
      col_done_2901 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2629_inst
    process(num_2611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_2611, konst_2628_wire_constant, tmp_var);
      EQ_u2_u1_2629_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2893_inst
    process(num_2611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_2611, konst_2892_wire_constant, tmp_var);
      EQ_u2_u1_2893_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2828_inst
    process(kval1_2816, ival1_2740) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_2816, ival1_2740, tmp_var);
      MUL_i16_i16_2828_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2834_inst
    process(kval2_2820, ival2_2744) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_2820, ival2_2744, tmp_var);
      MUL_i16_i16_2834_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2840_inst
    process(kval3_2824, ival3_2748) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_2824, ival3_2748, tmp_var);
      MUL_i16_i16_2840_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2846_inst
    process(kval1_2816, ival2_2744) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_2816, ival2_2744, tmp_var);
      MUL_i16_i16_2846_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2852_inst
    process(kval2_2820, ival3_2748) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_2820, ival3_2748, tmp_var);
      MUL_i16_i16_2852_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2858_inst
    process(kval3_2824, ival4_2752) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_2824, ival4_2752, tmp_var);
      MUL_i16_i16_2858_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2921_inst
    process(AND_u1_u1_2920_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AND_u1_u1_2920_wire, tmp_var);
      store_kernel_2922 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3023_inst
    process(all_done_flag_2927) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", all_done_flag_2927, tmp_var);
      NOT_u1_u1_3023_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2630_inst
    process(EQ_u16_u1_2626_wire, EQ_u2_u1_2629_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u16_u1_2626_wire, EQ_u2_u1_2629_wire, tmp_var);
      read_ip_2631 <= tmp_var; --
    end process;
    -- shared split operator group (32) : SUB_u16_u16_2576_inst 
    ApIntSub_group_32: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_2574_wire;
      num_row_2577 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2576_inst_req_0;
      SUB_u16_u16_2576_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2576_inst_req_1;
      SUB_u16_u16_2576_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_32_gI: SplitGuardInterface generic map(name => "ApIntSub_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : SUB_u16_u16_2581_inst 
    ApIntSub_group_33: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_2579_wire;
      num_col_2582 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2581_inst_req_0;
      SUB_u16_u16_2581_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2581_inst_req_1;
      SUB_u16_u16_2581_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_33_gI: SplitGuardInterface generic map(name => "ApIntSub_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : SUB_u16_u16_2586_inst 
    ApIntSub_group_34: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_size_pipe_2584_wire;
      num_chl_2587 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2586_inst_req_0;
      SUB_u16_u16_2586_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2586_inst_req_1;
      SUB_u16_u16_2586_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_34_gI: SplitGuardInterface generic map(name => "ApIntSub_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : SUB_u16_u16_2910_inst 
    ApIntSub_group_35: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= num_row_2577;
      SUB_u16_u16_2815_2815_delayed_1_0_2911 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2910_inst_req_0;
      SUB_u16_u16_2910_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2910_inst_req_1;
      SUB_u16_u16_2910_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_35_gI: SplitGuardInterface generic map(name => "ApIntSub_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- binary operator UGE_u16_u1_2915_inst
    process(row_2601, SUB_u16_u16_2815_2815_delayed_1_0_2911) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(row_2601, SUB_u16_u16_2815_2815_delayed_1_0_2911, tmp_var);
      out_done_flag_2916 <= tmp_var; --
    end process;
    -- binary operator UGT_u2_u1_2706_inst
    process(num_2611) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_2611, konst_2705_wire_constant, tmp_var);
      UGT_u2_u1_2706_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_2703_inst
    process(col_2606, num_col_2582) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(col_2606, num_col_2582, tmp_var);
      ULT_u16_u1_2703_wire <= tmp_var; --
    end process;
    xxconvolvexxconv_ip1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip1",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip1_pipe_read_req,
        read_ack => xxconvolvexxconv_ip1_pipe_read_ack,
        read_data => xxconvolvexxconv_ip1_pipe_read_data,
        write_req => xxconvolvexxconv_ip1_pipe_write_req,
        write_ack => xxconvolvexxconv_ip1_pipe_write_ack,
        write_data => xxconvolvexxconv_ip1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip2",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip2_pipe_read_req,
        read_ack => xxconvolvexxconv_ip2_pipe_read_ack,
        read_data => xxconvolvexxconv_ip2_pipe_read_data,
        write_req => xxconvolvexxconv_ip2_pipe_write_req,
        write_ack => xxconvolvexxconv_ip2_pipe_write_ack,
        write_data => xxconvolvexxconv_ip2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip3",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip3_pipe_read_req,
        read_ack => xxconvolvexxconv_ip3_pipe_read_ack,
        read_data => xxconvolvexxconv_ip3_pipe_read_data,
        write_req => xxconvolvexxconv_ip3_pipe_write_req,
        write_ack => xxconvolvexxconv_ip3_pipe_write_ack,
        write_data => xxconvolvexxconv_ip3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip4_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip4",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip4_pipe_read_req,
        read_ack => xxconvolvexxconv_ip4_pipe_read_ack,
        read_data => xxconvolvexxconv_ip4_pipe_read_data,
        write_req => xxconvolvexxconv_ip4_pipe_write_req,
        write_ack => xxconvolvexxconv_ip4_pipe_write_ack,
        write_data => xxconvolvexxconv_ip4_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k1",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k1_pipe_read_req,
        read_ack => xxconvolvexxconv_k1_pipe_read_ack,
        read_data => xxconvolvexxconv_k1_pipe_read_data,
        write_req => xxconvolvexxconv_k1_pipe_write_req,
        write_ack => xxconvolvexxconv_k1_pipe_write_ack,
        write_data => xxconvolvexxconv_k1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k2",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k2_pipe_read_req,
        read_ack => xxconvolvexxconv_k2_pipe_read_ack,
        read_data => xxconvolvexxconv_k2_pipe_read_data,
        write_req => xxconvolvexxconv_k2_pipe_write_req,
        write_ack => xxconvolvexxconv_k2_pipe_write_ack,
        write_data => xxconvolvexxconv_k2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k3",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k3_pipe_read_req,
        read_ack => xxconvolvexxconv_k3_pipe_read_ack,
        read_data => xxconvolvexxconv_k3_pipe_read_data,
        write_req => xxconvolvexxconv_k3_pipe_write_req,
        write_ack => xxconvolvexxconv_k3_pipe_write_ack,
        write_data => xxconvolvexxconv_k3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : RPIPE_input_pipe1_2634_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_2634_inst_req_0;
      RPIPE_input_pipe1_2634_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_2634_inst_req_1;
      RPIPE_input_pipe1_2634_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2631(0);
      temp2_1_2635 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_input_pipe2_2638_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe2_2638_inst_req_0;
      RPIPE_input_pipe2_2638_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe2_2638_inst_req_1;
      RPIPE_input_pipe2_2638_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2631(0);
      temp2_2_2639 <= data_out(15 downto 0);
      input_pipe2_read_1_gI: SplitGuardInterface generic map(name => "input_pipe2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe2_read_1: InputPortRevised -- 
        generic map ( name => "input_pipe2_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe2_pipe_read_req(0),
          oack => input_pipe2_pipe_read_ack(0),
          odata => input_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_input_pipe3_2642_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe3_2642_inst_req_0;
      RPIPE_input_pipe3_2642_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe3_2642_inst_req_1;
      RPIPE_input_pipe3_2642_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2631(0);
      temp2_3_2643 <= data_out(15 downto 0);
      input_pipe3_read_2_gI: SplitGuardInterface generic map(name => "input_pipe3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe3_read_2: InputPortRevised -- 
        generic map ( name => "input_pipe3_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe3_pipe_read_req(0),
          oack => input_pipe3_pipe_read_ack(0),
          odata => input_pipe3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_input_pipe4_2646_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe4_2646_inst_req_0;
      RPIPE_input_pipe4_2646_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe4_2646_inst_req_1;
      RPIPE_input_pipe4_2646_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_2631(0);
      temp2_4_2647 <= data_out(15 downto 0);
      input_pipe4_read_3_gI: SplitGuardInterface generic map(name => "input_pipe4_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe4_read_3: InputPortRevised -- 
        generic map ( name => "input_pipe4_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe4_pipe_read_req(0),
          oack => input_pipe4_pipe_read_ack(0),
          odata => input_pipe4_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_kernel_pipe1_2764_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_2764_inst_req_0;
      RPIPE_kernel_pipe1_2764_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_2764_inst_req_1;
      RPIPE_kernel_pipe1_2764_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2761(0);
      tempk1_1_2765 <= data_out(15 downto 0);
      kernel_pipe1_read_4_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_4: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_4", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : RPIPE_kernel_pipe2_2768_inst 
    InportGroup_5: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe2_2768_inst_req_0;
      RPIPE_kernel_pipe2_2768_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe2_2768_inst_req_1;
      RPIPE_kernel_pipe2_2768_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2761(0);
      tempk1_2_2769 <= data_out(15 downto 0);
      kernel_pipe2_read_5_gI: SplitGuardInterface generic map(name => "kernel_pipe2_read_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_read_5: InputPortRevised -- 
        generic map ( name => "kernel_pipe2_read_5", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe2_pipe_read_req(0),
          oack => kernel_pipe2_pipe_read_ack(0),
          odata => kernel_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : RPIPE_kernel_pipe3_2772_inst 
    InportGroup_6: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe3_2772_inst_req_0;
      RPIPE_kernel_pipe3_2772_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe3_2772_inst_req_1;
      RPIPE_kernel_pipe3_2772_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2761(0);
      tempk1_3_2773 <= data_out(15 downto 0);
      kernel_pipe3_read_6_gI: SplitGuardInterface generic map(name => "kernel_pipe3_read_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_read_6: InputPortRevised -- 
        generic map ( name => "kernel_pipe3_read_6", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe3_pipe_read_req(0),
          oack => kernel_pipe3_pipe_read_ack(0),
          odata => kernel_pipe3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : RPIPE_num_out_pipe_2574_inst RPIPE_num_out_pipe_2579_inst 
    InportGroup_7: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_num_out_pipe_2574_inst_req_0;
      reqL_unguarded(0) <= RPIPE_num_out_pipe_2579_inst_req_0;
      RPIPE_num_out_pipe_2574_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_num_out_pipe_2579_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_num_out_pipe_2574_inst_req_1;
      reqR_unguarded(0) <= RPIPE_num_out_pipe_2579_inst_req_1;
      RPIPE_num_out_pipe_2574_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_num_out_pipe_2579_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      RPIPE_num_out_pipe_2574_wire <= data_out(31 downto 16);
      RPIPE_num_out_pipe_2579_wire <= data_out(15 downto 0);
      num_out_pipe_read_7_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_7_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_7: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_7", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : RPIPE_size_pipe_2584_inst 
    InportGroup_8: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_2584_inst_req_0;
      RPIPE_size_pipe_2584_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_2584_inst_req_1;
      RPIPE_size_pipe_2584_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_size_pipe_2584_wire <= data_out(15 downto 0);
      size_pipe_read_8_gI: SplitGuardInterface generic map(name => "size_pipe_read_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_8: InputPortRevised -- 
        generic map ( name => "size_pipe_read_8", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : RPIPE_xxconvolvexxconv_ip1_2650_inst 
    InportGroup_9: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_2650_inst_req_0;
      RPIPE_xxconvolvexxconv_ip1_2650_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_2650_inst_req_1;
      RPIPE_xxconvolvexxconv_ip1_2650_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2631(0);
      temp1_1_2651 <= data_out(15 downto 0);
      xxconvolvexxconv_ip1_read_9_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_read_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_read_9: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1_read_9", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip1_pipe_read_req(0),
          oack => xxconvolvexxconv_ip1_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : RPIPE_xxconvolvexxconv_ip2_2654_inst 
    InportGroup_10: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_2654_inst_req_0;
      RPIPE_xxconvolvexxconv_ip2_2654_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_2654_inst_req_1;
      RPIPE_xxconvolvexxconv_ip2_2654_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2631(0);
      temp1_2_2655 <= data_out(15 downto 0);
      xxconvolvexxconv_ip2_read_10_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_read_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_read_10: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2_read_10", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip2_pipe_read_req(0),
          oack => xxconvolvexxconv_ip2_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : RPIPE_xxconvolvexxconv_ip3_2658_inst 
    InportGroup_11: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_2658_inst_req_0;
      RPIPE_xxconvolvexxconv_ip3_2658_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_2658_inst_req_1;
      RPIPE_xxconvolvexxconv_ip3_2658_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2631(0);
      temp1_3_2659 <= data_out(15 downto 0);
      xxconvolvexxconv_ip3_read_11_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_read_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_read_11: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3_read_11", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip3_pipe_read_req(0),
          oack => xxconvolvexxconv_ip3_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- shared inport operator group (12) : RPIPE_xxconvolvexxconv_ip4_2662_inst 
    InportGroup_12: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip4_2662_inst_req_0;
      RPIPE_xxconvolvexxconv_ip4_2662_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip4_2662_inst_req_1;
      RPIPE_xxconvolvexxconv_ip4_2662_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_2631(0);
      temp1_4_2663 <= data_out(15 downto 0);
      xxconvolvexxconv_ip4_read_12_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip4_read_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip4_read_12: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip4_read_12", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip4_pipe_read_req(0),
          oack => xxconvolvexxconv_ip4_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip4_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 12
    -- shared inport operator group (13) : RPIPE_xxconvolvexxconv_k1_2776_inst 
    InportGroup_13: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2776_inst_req_0;
      RPIPE_xxconvolvexxconv_k1_2776_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2776_inst_req_1;
      RPIPE_xxconvolvexxconv_k1_2776_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2761(0);
      tempk2_1_2777 <= data_out(15 downto 0);
      xxconvolvexxconv_k1_read_13_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_read_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_read_13: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1_read_13", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k1_pipe_read_req(0),
          oack => xxconvolvexxconv_k1_pipe_read_ack(0),
          odata => xxconvolvexxconv_k1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 13
    -- shared inport operator group (14) : RPIPE_xxconvolvexxconv_k2_2780_inst 
    InportGroup_14: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2780_inst_req_0;
      RPIPE_xxconvolvexxconv_k2_2780_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2780_inst_req_1;
      RPIPE_xxconvolvexxconv_k2_2780_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2761(0);
      tempk2_2_2781 <= data_out(15 downto 0);
      xxconvolvexxconv_k2_read_14_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_read_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_read_14: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2_read_14", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k2_pipe_read_req(0),
          oack => xxconvolvexxconv_k2_pipe_read_ack(0),
          odata => xxconvolvexxconv_k2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 14
    -- shared inport operator group (15) : RPIPE_xxconvolvexxconv_k3_2784_inst 
    InportGroup_15: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2784_inst_req_0;
      RPIPE_xxconvolvexxconv_k3_2784_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2784_inst_req_1;
      RPIPE_xxconvolvexxconv_k3_2784_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2761(0);
      tempk2_3_2785 <= data_out(15 downto 0);
      xxconvolvexxconv_k3_read_15_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_read_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_read_15: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3_read_15", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k3_pipe_read_req(0),
          oack => xxconvolvexxconv_k3_pipe_read_ack(0),
          odata => xxconvolvexxconv_k3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 15
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3024_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3024_inst_req_0;
      WPIPE_input_done_pipe_3024_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3024_inst_req_1;
      WPIPE_input_done_pipe_3024_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3025_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_output_pipe_3009_inst WPIPE_output_pipe_3017_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_output_pipe_3009_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_output_pipe_3017_inst_req_0;
      WPIPE_output_pipe_3009_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_output_pipe_3017_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_output_pipe_3009_inst_req_1;
      update_req_unguarded(0) <= WPIPE_output_pipe_3017_inst_req_1;
      WPIPE_output_pipe_3009_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_output_pipe_3017_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= num_done_2896_delayed_1_0_3015(0);
      guard_vector(1)  <= num_done_2891_delayed_1_0_3007(0);
      data_in <= type_cast_3011_wire & type_cast_3019_wire;
      output_pipe_write_1_gI: SplitGuardInterface generic map(name => "output_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_xxconvolvexxconv_ip1_2713_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2713_inst_req_0;
      WPIPE_xxconvolvexxconv_ip1_2713_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2713_inst_req_1;
      WPIPE_xxconvolvexxconv_ip1_2713_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2640_delayed_1_0_2711(0);
      data_in <= iread1_2672;
      xxconvolvexxconv_ip1_write_2_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_write_2: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip1_pipe_write_req(0),
          oack => xxconvolvexxconv_ip1_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_xxconvolvexxconv_ip2_2720_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2720_inst_req_0;
      WPIPE_xxconvolvexxconv_ip2_2720_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2720_inst_req_1;
      WPIPE_xxconvolvexxconv_ip2_2720_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2644_delayed_1_0_2718(0);
      data_in <= iread2_2681;
      xxconvolvexxconv_ip2_write_3_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_write_3: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip2_pipe_write_req(0),
          oack => xxconvolvexxconv_ip2_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_xxconvolvexxconv_ip3_2727_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2727_inst_req_0;
      WPIPE_xxconvolvexxconv_ip3_2727_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2727_inst_req_1;
      WPIPE_xxconvolvexxconv_ip3_2727_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2648_delayed_1_0_2725(0);
      data_in <= iread3_2690;
      xxconvolvexxconv_ip3_write_4_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_write_4: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip3_pipe_write_req(0),
          oack => xxconvolvexxconv_ip3_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_xxconvolvexxconv_ip4_2734_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip4_2734_inst_req_0;
      WPIPE_xxconvolvexxconv_ip4_2734_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip4_2734_inst_req_1;
      WPIPE_xxconvolvexxconv_ip4_2734_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_2652_delayed_1_0_2732(0);
      data_in <= iread4_2699;
      xxconvolvexxconv_ip4_write_5_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip4_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip4_write_5: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip4", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip4_pipe_write_req(0),
          oack => xxconvolvexxconv_ip4_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip4_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_xxconvolvexxconv_k1_2932_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_2932_inst_req_0;
      WPIPE_xxconvolvexxconv_k1_2932_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_2932_inst_req_1;
      WPIPE_xxconvolvexxconv_k1_2932_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2829_delayed_1_0_2930(0);
      data_in <= kread1_2794;
      xxconvolvexxconv_k1_write_6_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_write_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_write_6: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k1_pipe_write_req(0),
          oack => xxconvolvexxconv_k1_pipe_write_ack(0),
          odata => xxconvolvexxconv_k1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_xxconvolvexxconv_k2_2939_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_2939_inst_req_0;
      WPIPE_xxconvolvexxconv_k2_2939_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_2939_inst_req_1;
      WPIPE_xxconvolvexxconv_k2_2939_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2833_delayed_1_0_2937(0);
      data_in <= kread2_2803;
      xxconvolvexxconv_k2_write_7_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_write_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_write_7: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k2_pipe_write_req(0),
          oack => xxconvolvexxconv_k2_pipe_write_ack(0),
          odata => xxconvolvexxconv_k2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- shared outport operator group (8) : WPIPE_xxconvolvexxconv_k3_2946_inst 
    OutportGroup_8: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_2946_inst_req_0;
      WPIPE_xxconvolvexxconv_k3_2946_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_2946_inst_req_1;
      WPIPE_xxconvolvexxconv_k3_2946_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2837_delayed_1_0_2944(0);
      data_in <= kread3_2812;
      xxconvolvexxconv_k3_write_8_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_write_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_write_8: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k3_pipe_write_req(0),
          oack => xxconvolvexxconv_k3_pipe_write_ack(0),
          odata => xxconvolvexxconv_k3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    num_chl : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal num_chl_buffer :  std_logic_vector(15 downto 0);
  signal num_chl_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_1635_start: Boolean;
  signal loadKernelChannel_CP_1635_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_kernel_pipe1_629_inst_ack_0 : boolean;
  signal addr_of_543_final_reg_ack_1 : boolean;
  signal array_obj_ref_542_index_offset_ack_0 : boolean;
  signal phi_stmt_581_req_0 : boolean;
  signal start_add_583_buf_ack_0 : boolean;
  signal addr_of_543_final_reg_req_1 : boolean;
  signal my_fetch_548_587_buf_req_1 : boolean;
  signal do_while_stmt_579_branch_req_0 : boolean;
  signal phi_stmt_585_req_1 : boolean;
  signal addr_of_543_final_reg_ack_0 : boolean;
  signal array_obj_ref_542_index_offset_req_0 : boolean;
  signal phi_stmt_581_req_1 : boolean;
  signal RPIPE_input_done_pipe_576_inst_req_0 : boolean;
  signal array_obj_ref_542_index_offset_ack_1 : boolean;
  signal ptr_deref_547_load_0_req_0 : boolean;
  signal RPIPE_input_done_pipe_576_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_576_inst_req_1 : boolean;
  signal ptr_deref_547_load_0_ack_0 : boolean;
  signal ptr_deref_547_load_0_req_1 : boolean;
  signal RPIPE_input_done_pipe_576_inst_ack_0 : boolean;
  signal phi_stmt_581_ack_0 : boolean;
  signal addr_of_543_final_reg_req_0 : boolean;
  signal my_fetch_548_587_buf_req_0 : boolean;
  signal nmycount_603_584_buf_ack_0 : boolean;
  signal nmycount_603_584_buf_req_0 : boolean;
  signal start_add_583_buf_ack_1 : boolean;
  signal ptr_deref_547_load_0_ack_1 : boolean;
  signal nmycount_603_584_buf_ack_1 : boolean;
  signal nmycount_603_584_buf_req_1 : boolean;
  signal phi_stmt_585_req_0 : boolean;
  signal my_fetch_548_587_buf_ack_1 : boolean;
  signal nfetch_val_675_588_buf_req_1 : boolean;
  signal nfetch_val_675_588_buf_ack_0 : boolean;
  signal array_obj_ref_542_index_offset_req_1 : boolean;
  signal WPIPE_kernel_pipe1_629_inst_ack_1 : boolean;
  signal nfetch_val_675_588_buf_req_0 : boolean;
  signal phi_stmt_585_ack_0 : boolean;
  signal start_add_583_buf_req_0 : boolean;
  signal WPIPE_kernel_pipe1_629_inst_req_1 : boolean;
  signal array_obj_ref_653_index_offset_req_0 : boolean;
  signal array_obj_ref_653_index_offset_ack_0 : boolean;
  signal start_add_583_buf_req_1 : boolean;
  signal WPIPE_kernel_pipe2_633_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_633_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe3_637_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe3_637_inst_ack_1 : boolean;
  signal array_obj_ref_653_index_offset_req_1 : boolean;
  signal array_obj_ref_653_index_offset_ack_1 : boolean;
  signal addr_of_654_final_reg_req_0 : boolean;
  signal WPIPE_kernel_pipe1_629_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_633_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_633_inst_ack_1 : boolean;
  signal my_fetch_548_587_buf_ack_0 : boolean;
  signal WPIPE_kernel_pipe3_637_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe3_637_inst_ack_0 : boolean;
  signal nfetch_val_675_588_buf_ack_1 : boolean;
  signal addr_of_654_final_reg_ack_0 : boolean;
  signal addr_of_654_final_reg_req_1 : boolean;
  signal addr_of_654_final_reg_ack_1 : boolean;
  signal W_fn_608_delayed_7_0_656_inst_req_0 : boolean;
  signal W_fn_608_delayed_7_0_656_inst_ack_0 : boolean;
  signal W_fn_608_delayed_7_0_656_inst_req_1 : boolean;
  signal W_fn_608_delayed_7_0_656_inst_ack_1 : boolean;
  signal ptr_deref_662_load_0_req_0 : boolean;
  signal ptr_deref_662_load_0_ack_0 : boolean;
  signal ptr_deref_662_load_0_req_1 : boolean;
  signal ptr_deref_662_load_0_ack_1 : boolean;
  signal W_fn_614_delayed_13_0_664_inst_req_0 : boolean;
  signal W_fn_614_delayed_13_0_664_inst_ack_0 : boolean;
  signal W_fn_614_delayed_13_0_664_inst_req_1 : boolean;
  signal W_fn_614_delayed_13_0_664_inst_ack_1 : boolean;
  signal W_fetch_val_616_delayed_13_0_667_inst_req_0 : boolean;
  signal W_fetch_val_616_delayed_13_0_667_inst_ack_0 : boolean;
  signal W_fetch_val_616_delayed_13_0_667_inst_req_1 : boolean;
  signal W_fetch_val_616_delayed_13_0_667_inst_ack_1 : boolean;
  signal do_while_stmt_579_branch_ack_0 : boolean;
  signal do_while_stmt_579_branch_ack_1 : boolean;
  signal WPIPE_size_pipe_683_inst_req_0 : boolean;
  signal WPIPE_size_pipe_683_inst_ack_0 : boolean;
  signal WPIPE_size_pipe_683_inst_req_1 : boolean;
  signal WPIPE_size_pipe_683_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(79 downto 64) <= num_chl;
  num_chl_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_1635_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1635_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1635_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1635_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_1635: Block -- control-path 
    signal loadKernelChannel_CP_1635_elements: BooleanArray(98 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_1635_elements(0) <= loadKernelChannel_CP_1635_start;
    loadKernelChannel_CP_1635_symbol <= loadKernelChannel_CP_1635_elements(98);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_complete/req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_update_start_
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_sample_start_
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Sample/rr
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_complete/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_computed_1
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_index_resized_1
      -- CP-element group 0: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_update_start_
      -- 
    req_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => array_obj_ref_542_index_offset_req_0); -- 
    req_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => array_obj_ref_542_index_offset_req_1); -- 
    req_1685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => addr_of_543_final_reg_req_1); -- 
    cr_1730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => ptr_deref_547_load_0_req_1); -- 
    rr_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(0), ack => RPIPE_input_done_pipe_576_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Sample/ack
      -- CP-element group 1: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_sample_complete
      -- 
    ack_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_542_index_offset_ack_0, ack => loadKernelChannel_CP_1635_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_request/req
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_request/$entry
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_sample_start_
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_offset_calculated
      -- CP-element group 2: 	 assign_stmt_532_to_assign_stmt_577/array_obj_ref_542_root_address_calculated
      -- 
    ack_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_542_index_offset_ack_1, ack => loadKernelChannel_CP_1635_elements(2)); -- 
    req_1680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(2), ack => addr_of_543_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_sample_completed_
      -- CP-element group 3: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_request/ack
      -- CP-element group 3: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_request/$exit
      -- 
    ack_1681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_543_final_reg_ack_0, ack => loadKernelChannel_CP_1635_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_complete/ack
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_sample_start_
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_address_resized
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/word_0/rr
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_complete/$exit
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_532_to_assign_stmt_577/addr_of_543_update_completed_
      -- 
    ack_1686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_543_final_reg_ack_1, ack => loadKernelChannel_CP_1635_elements(4)); -- 
    rr_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(4), ack => ptr_deref_547_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_sample_completed_
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Sample/$exit
      -- 
    ra_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_547_load_0_ack_0, ack => loadKernelChannel_CP_1635_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/ptr_deref_547_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/ptr_deref_547_Merge/merge_ack
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_update_completed_
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/ptr_deref_547_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/ptr_deref_547_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/$exit
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_532_to_assign_stmt_577/ptr_deref_547_Update/word_access_complete/word_0/$exit
      -- 
    ca_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_547_load_0_ack_1, ack => loadKernelChannel_CP_1635_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Update/cr
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Update/$entry
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Sample/ra
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_update_start_
      -- CP-element group 7: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_sample_completed_
      -- 
    ra_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_576_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(7)); -- 
    cr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(7), ack => RPIPE_input_done_pipe_576_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Update/ca
      -- CP-element group 8: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_Update/$exit
      -- CP-element group 8: 	 assign_stmt_532_to_assign_stmt_577/RPIPE_input_done_pipe_576_update_completed_
      -- 
    ca_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_576_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_578/branch_block_stmt_578__entry__
      -- CP-element group 9: 	 branch_block_stmt_578/$entry
      -- CP-element group 9: 	 branch_block_stmt_578/do_while_stmt_579__entry__
      -- CP-element group 9: 	 assign_stmt_532_to_assign_stmt_577/$exit
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(1) & loadKernelChannel_CP_1635_elements(6) & loadKernelChannel_CP_1635_elements(8);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	96 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	97 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_578/$exit
      -- CP-element group 10: 	 branch_block_stmt_578/branch_block_stmt_578__exit__
      -- CP-element group 10: 	 branch_block_stmt_578/do_while_stmt_579__exit__
      -- CP-element group 10: 	 assign_stmt_685/$entry
      -- CP-element group 10: 	 assign_stmt_685/WPIPE_size_pipe_683_sample_start_
      -- CP-element group 10: 	 assign_stmt_685/WPIPE_size_pipe_683_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_685/WPIPE_size_pipe_683_Sample/req
      -- 
    req_2086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(10), ack => WPIPE_size_pipe_683_inst_req_0); -- 
    loadKernelChannel_CP_1635_elements(10) <= loadKernelChannel_CP_1635_elements(96);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_578/do_while_stmt_579/$entry
      -- CP-element group 11: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579__entry__
      -- 
    loadKernelChannel_CP_1635_elements(11) <= loadKernelChannel_CP_1635_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	96 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579__exit__
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_578/do_while_stmt_579/loop_back
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	94 
    -- CP-element group 14: 	95 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_578/do_while_stmt_579/condition_done
      -- CP-element group 14: 	 branch_block_stmt_578/do_while_stmt_579/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_578/do_while_stmt_579/loop_taken/$entry
      -- 
    loadKernelChannel_CP_1635_elements(14) <= loadKernelChannel_CP_1635_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	93 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_578/do_while_stmt_579/loop_body_done
      -- 
    loadKernelChannel_CP_1635_elements(15) <= loadKernelChannel_CP_1635_elements(93);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	28 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_1635_elements(16) <= loadKernelChannel_CP_1635_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_1635_elements(17) <= loadKernelChannel_CP_1635_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	70 
    -- CP-element group 18: 	71 
    -- CP-element group 18: 	92 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	27 
    -- CP-element group 19: 	92 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/condition_evaluated
      -- 
    condition_evaluated_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(19), ack => do_while_stmt_579_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(23) & loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(92);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	41 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/aggregated_phi_sample_req
      -- CP-element group 20: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_sample_start__ps
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(24) & loadKernelChannel_CP_1635_elements(41) & loadKernelChannel_CP_1635_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	81 
    -- CP-element group 21: 	85 
    -- CP-element group 21: 	89 
    -- CP-element group 21: 	93 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	41 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(26) & loadKernelChannel_CP_1635_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	42 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/aggregated_phi_update_req
      -- CP-element group 22: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_update_start__ps
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(25) & loadKernelChannel_CP_1635_elements(42);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	64 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	78 
    -- CP-element group 25: 	86 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(61) & loadKernelChannel_CP_1635_elements(64) & loadKernelChannel_CP_1635_elements(67) & loadKernelChannel_CP_1635_elements(72) & loadKernelChannel_CP_1635_elements(78) & loadKernelChannel_CP_1635_elements(86);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	23 
    -- CP-element group 27: 	60 
    -- CP-element group 27: 	63 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	72 
    -- CP-element group 27: 	76 
    -- CP-element group 27: 	84 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (15) 
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_index_resize_1/index_resize_ack
      -- 
    req_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(27), ack => array_obj_ref_653_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	16 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_loopback_trigger
      -- 
    loadKernelChannel_CP_1635_elements(28) <= loadKernelChannel_CP_1635_elements(16);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_loopback_sample_req
      -- CP-element group 29: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_loopback_sample_req_ps
      -- 
    phi_stmt_581_loopback_sample_req_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_581_loopback_sample_req_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(29), ack => phi_stmt_581_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_entry_trigger
      -- 
    loadKernelChannel_CP_1635_elements(30) <= loadKernelChannel_CP_1635_elements(17);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_entry_sample_req
      -- CP-element group 31: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_entry_sample_req_ps
      -- 
    phi_stmt_581_entry_sample_req_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_581_entry_sample_req_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(31), ack => phi_stmt_581_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_phi_mux_ack_ps
      -- CP-element group 32: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_581_phi_mux_ack
      -- 
    phi_stmt_581_phi_mux_ack_1793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_581_ack_0, ack => loadKernelChannel_CP_1635_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Sample/req
      -- 
    req_1806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(33), ack => start_add_583_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_update_start_
      -- CP-element group 34: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Update/req
      -- CP-element group 34: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Update/$entry
      -- 
    req_1811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(34), ack => start_add_583_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Sample/ack
      -- CP-element group 35: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Sample/$exit
      -- 
    ack_1807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_583_buf_ack_0, ack => loadKernelChannel_CP_1635_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_start_add_583_Update/$exit
      -- 
    ack_1812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_583_buf_ack_1, ack => loadKernelChannel_CP_1635_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_sample_start__ps
      -- CP-element group 37: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Sample/$entry
      -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(37), ack => nmycount_603_584_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Update/req
      -- CP-element group 38: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_update_start_
      -- 
    req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(38), ack => nmycount_603_584_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Sample/$exit
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_603_584_buf_ack_0, ack => loadKernelChannel_CP_1635_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nmycount_584_update_completed_
      -- 
    ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_603_584_buf_ack_1, ack => loadKernelChannel_CP_1635_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	21 
    -- CP-element group 41: 	83 
    -- CP-element group 41: 	87 
    -- CP-element group 41: 	91 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_sample_start_
      -- 
    loadKernelChannel_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(83) & loadKernelChannel_CP_1635_elements(87) & loadKernelChannel_CP_1635_elements(91);
      gj_loadKernelChannel_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	46 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	64 
    -- CP-element group 42: 	67 
    -- CP-element group 42: 	90 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	22 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_update_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(61) & loadKernelChannel_CP_1635_elements(64) & loadKernelChannel_CP_1635_elements(67) & loadKernelChannel_CP_1635_elements(90);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_sample_start__ps
      -- 
    loadKernelChannel_CP_1635_elements(43) <= loadKernelChannel_CP_1635_elements(20);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_update_start__ps
      -- 
    loadKernelChannel_CP_1635_elements(45) <= loadKernelChannel_CP_1635_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	63 
    -- CP-element group 46: 	66 
    -- CP-element group 46: 	88 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_update_completed_
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_loopback_trigger
      -- 
    loadKernelChannel_CP_1635_elements(47) <= loadKernelChannel_CP_1635_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_loopback_sample_req
      -- CP-element group 48: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_loopback_sample_req_ps
      -- 
    phi_stmt_585_loopback_sample_req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_585_loopback_sample_req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(48), ack => phi_stmt_585_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_entry_trigger
      -- 
    loadKernelChannel_CP_1635_elements(49) <= loadKernelChannel_CP_1635_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_entry_sample_req_ps
      -- CP-element group 50: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_entry_sample_req
      -- 
    phi_stmt_585_entry_sample_req_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_585_entry_sample_req_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(50), ack => phi_stmt_585_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/phi_stmt_585_phi_mux_ack_ps
      -- 
    phi_stmt_585_phi_mux_ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_585_ack_0, ack => loadKernelChannel_CP_1635_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_Sample/$entry
      -- 
    req_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(52), ack => my_fetch_548_587_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_Update/req
      -- CP-element group 53: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_update_start_
      -- 
    req_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(53), ack => my_fetch_548_587_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_Sample/ack
      -- 
    ack_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_548_587_buf_ack_0, ack => loadKernelChannel_CP_1635_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_my_fetch_587_Update/ack
      -- 
    ack_1866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_548_587_buf_ack_1, ack => loadKernelChannel_CP_1635_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_Sample/req
      -- 
    req_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(56), ack => nfetch_val_675_588_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1635_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_update_start_
      -- CP-element group 57: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_Update/req
      -- CP-element group 57: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_update_start__ps
      -- 
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(57), ack => nfetch_val_675_588_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1635_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_sample_completed__ps
      -- 
    ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_675_588_buf_ack_0, ack => loadKernelChannel_CP_1635_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_update_completed__ps
      -- CP-element group 59: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/R_nfetch_val_588_Update/ack
      -- 
    ack_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_675_588_buf_ack_1, ack => loadKernelChannel_CP_1635_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Sample/req
      -- 
    req_1893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(60), ack => WPIPE_kernel_pipe1_629_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	25 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_update_start_
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Update/req
      -- 
    ack_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_629_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(61)); -- 
    req_1898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(61), ack => WPIPE_kernel_pipe1_629_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	93 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe1_629_update_completed_
      -- 
    ack_1899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_629_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	27 
    -- CP-element group 63: 	46 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_sample_start_
      -- 
    req_1907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(63), ack => WPIPE_kernel_pipe2_633_inst_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(65);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	25 
    -- CP-element group 64: 	42 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Update/req
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_update_start_
      -- 
    ack_1908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_633_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(64)); -- 
    req_1912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(64), ack => WPIPE_kernel_pipe2_633_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	93 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe2_633_Update/ack
      -- 
    ack_1913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_633_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	27 
    -- CP-element group 66: 	46 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Sample/req
      -- 
    req_1921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(66), ack => WPIPE_kernel_pipe3_637_inst_req_0); -- 
    loadKernelChannel_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(68);
      gj_loadKernelChannel_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	42 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_update_start_
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Update/req
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Update/$entry
      -- 
    ack_1922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_637_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(67)); -- 
    req_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(67), ack => WPIPE_kernel_pipe3_637_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	93 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/WPIPE_kernel_pipe3_637_update_completed_
      -- 
    ack_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_637_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	73 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_request/$entry
      -- CP-element group 69: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_request/req
      -- CP-element group 69: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_sample_start_
      -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(69), ack => addr_of_654_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(73) & loadKernelChannel_CP_1635_elements(74);
      gj_loadKernelChannel_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	18 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	75 
    -- CP-element group 70: 	82 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	75 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_update_start_
      -- CP-element group 70: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_complete/$entry
      -- CP-element group 70: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_complete/req
      -- 
    req_1972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(70), ack => addr_of_654_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(75) & loadKernelChannel_CP_1635_elements(82);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	18 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	74 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_update_start
      -- CP-element group 71: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Update/req
      -- 
    req_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(71), ack => array_obj_ref_653_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(18) & loadKernelChannel_CP_1635_elements(73) & loadKernelChannel_CP_1635_elements(74);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	27 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	93 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_sample_complete
      -- CP-element group 72: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Sample/ack
      -- 
    ack_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_653_index_offset_ack_0, ack => loadKernelChannel_CP_1635_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (8) 
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_offset_calculated
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_final_index_sum_regn_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/array_obj_ref_653_base_plus_offset/sum_rename_ack
      -- 
    ack_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_653_index_offset_ack_1, ack => loadKernelChannel_CP_1635_elements(73)); -- 
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	71 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_request/$exit
      -- CP-element group 74: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_request/ack
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_654_final_reg_ack_0, ack => loadKernelChannel_CP_1635_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	70 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	80 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	70 
    -- CP-element group 75:  members (19) 
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/addr_of_654_complete/ack
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_root_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_address_resized
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_addr_resize/$entry
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_addr_resize/$exit
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_addr_resize/base_resize_req
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_addr_resize/base_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_plus_offset/$entry
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_plus_offset/$exit
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_plus_offset/sum_rename_req
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_base_plus_offset/sum_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_addrgen/$entry
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_addrgen/$exit
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_addrgen/root_register_req
      -- CP-element group 75: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_word_addrgen/root_register_ack
      -- 
    ack_1973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_654_final_reg_ack_1, ack => loadKernelChannel_CP_1635_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	27 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Sample/req
      -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(76), ack => W_fn_608_delayed_7_0_656_inst_req_0); -- 
    loadKernelChannel_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(78);
      gj_loadKernelChannel_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	82 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_update_start_
      -- CP-element group 77: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Update/req
      -- 
    req_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(77), ack => W_fn_608_delayed_7_0_656_inst_req_1); -- 
    loadKernelChannel_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(79) & loadKernelChannel_CP_1635_elements(82);
      gj_loadKernelChannel_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	25 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Sample/ack
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_608_delayed_7_0_656_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_658_Update/ack
      -- 
    ack_1987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_608_delayed_7_0_656_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: 	79 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/word_0/rr
      -- 
    rr_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(80), ack => ptr_deref_662_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(75) & loadKernelChannel_CP_1635_elements(79) & loadKernelChannel_CP_1635_elements(82);
      gj_loadKernelChannel_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	21 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_update_start_
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/word_0/cr
      -- 
    cr_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(81), ack => ptr_deref_662_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(83);
      gj_loadKernelChannel_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/$exit
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Sample/word_access_start/word_0/ra
      -- 
    ra_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_662_load_0_ack_0, ack => loadKernelChannel_CP_1635_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	93 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	41 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/$exit
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/word_access_complete/word_0/ca
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/ptr_deref_662_Merge/$entry
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/ptr_deref_662_Merge/$exit
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/ptr_deref_662_Merge/merge_req
      -- CP-element group 83: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/ptr_deref_662_Update/ptr_deref_662_Merge/merge_ack
      -- 
    ca_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_662_load_0_ack_1, ack => loadKernelChannel_CP_1635_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	27 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Sample/req
      -- 
    req_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(84), ack => W_fn_614_delayed_13_0_664_inst_req_0); -- 
    loadKernelChannel_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(27) & loadKernelChannel_CP_1635_elements(86);
      gj_loadKernelChannel_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	21 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_update_start_
      -- CP-element group 85: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Update/req
      -- 
    req_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(85), ack => W_fn_614_delayed_13_0_664_inst_req_1); -- 
    loadKernelChannel_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(87);
      gj_loadKernelChannel_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	25 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Sample/ack
      -- 
    ack_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_614_delayed_13_0_664_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	93 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_666_Update/ack
      -- 
    ack_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_614_delayed_13_0_664_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	46 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Sample/req
      -- 
    req_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(88), ack => W_fetch_val_616_delayed_13_0_667_inst_req_0); -- 
    loadKernelChannel_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(46) & loadKernelChannel_CP_1635_elements(90);
      gj_loadKernelChannel_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	21 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_update_start_
      -- CP-element group 89: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Update/req
      -- 
    req_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(89), ack => W_fetch_val_616_delayed_13_0_667_inst_req_1); -- 
    loadKernelChannel_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(91);
      gj_loadKernelChannel_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	42 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Sample/ack
      -- 
    ack_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_616_delayed_13_0_667_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	41 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/assign_stmt_669_Update/ack
      -- 
    ack_2065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_616_delayed_13_0_667_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(91)); -- 
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	18 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	19 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_1635_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_1635_elements(18), ack => loadKernelChannel_CP_1635_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	21 
    -- CP-element group 93: 	62 
    -- CP-element group 93: 	65 
    -- CP-element group 93: 	68 
    -- CP-element group 93: 	72 
    -- CP-element group 93: 	83 
    -- CP-element group 93: 	87 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	15 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_578/do_while_stmt_579/do_while_stmt_579_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1635_elements(21) & loadKernelChannel_CP_1635_elements(62) & loadKernelChannel_CP_1635_elements(65) & loadKernelChannel_CP_1635_elements(68) & loadKernelChannel_CP_1635_elements(72) & loadKernelChannel_CP_1635_elements(83) & loadKernelChannel_CP_1635_elements(87) & loadKernelChannel_CP_1635_elements(91);
      gj_loadKernelChannel_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_578/do_while_stmt_579/loop_exit/$exit
      -- CP-element group 94: 	 branch_block_stmt_578/do_while_stmt_579/loop_exit/ack
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_579_branch_ack_0, ack => loadKernelChannel_CP_1635_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	14 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_578/do_while_stmt_579/loop_taken/$exit
      -- CP-element group 95: 	 branch_block_stmt_578/do_while_stmt_579/loop_taken/ack
      -- 
    ack_2074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_579_branch_ack_1, ack => loadKernelChannel_CP_1635_elements(95)); -- 
    -- CP-element group 96:  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	12 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	10 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_578/do_while_stmt_579/$exit
      -- 
    loadKernelChannel_CP_1635_elements(96) <= loadKernelChannel_CP_1635_elements(12);
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	10 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_sample_completed_
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_update_start_
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_Sample/$exit
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_Sample/ack
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_Update/$entry
      -- CP-element group 97: 	 assign_stmt_685/WPIPE_size_pipe_683_Update/req
      -- 
    ack_2087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_683_inst_ack_0, ack => loadKernelChannel_CP_1635_elements(97)); -- 
    req_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1635_elements(97), ack => WPIPE_size_pipe_683_inst_req_1); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 $exit
      -- CP-element group 98: 	 assign_stmt_685/$exit
      -- CP-element group 98: 	 assign_stmt_685/WPIPE_size_pipe_683_update_completed_
      -- CP-element group 98: 	 assign_stmt_685/WPIPE_size_pipe_683_Update/$exit
      -- CP-element group 98: 	 assign_stmt_685/WPIPE_size_pipe_683_Update/ack
      -- 
    ack_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_683_inst_ack_1, ack => loadKernelChannel_CP_1635_elements(98)); -- 
    loadKernelChannel_do_while_stmt_579_terminator_2075: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_579_terminator_2075", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_1635_elements(15),loop_continue => loadKernelChannel_CP_1635_elements(95),loop_terminate => loadKernelChannel_CP_1635_elements(94),loop_back => loadKernelChannel_CP_1635_elements(13),loop_exit => loadKernelChannel_CP_1635_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_581_phi_seq_1831_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1635_elements(30);
      loadKernelChannel_CP_1635_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1635_elements(35);
      loadKernelChannel_CP_1635_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1635_elements(36);
      loadKernelChannel_CP_1635_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1635_elements(28);
      loadKernelChannel_CP_1635_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1635_elements(39);
      loadKernelChannel_CP_1635_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1635_elements(40);
      loadKernelChannel_CP_1635_elements(29) <= phi_mux_reqs(1);
      phi_stmt_581_phi_seq_1831 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_581_phi_seq_1831") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1635_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_1635_elements(26), 
          phi_update_req => loadKernelChannel_CP_1635_elements(22), 
          phi_update_ack => loadKernelChannel_CP_1635_elements(27), 
          phi_mux_ack => loadKernelChannel_CP_1635_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_585_phi_seq_1885_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1635_elements(49);
      loadKernelChannel_CP_1635_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1635_elements(54);
      loadKernelChannel_CP_1635_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1635_elements(55);
      loadKernelChannel_CP_1635_elements(50) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1635_elements(47);
      loadKernelChannel_CP_1635_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1635_elements(58);
      loadKernelChannel_CP_1635_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1635_elements(59);
      loadKernelChannel_CP_1635_elements(48) <= phi_mux_reqs(1);
      phi_stmt_585_phi_seq_1885 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_585_phi_seq_1885") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1635_elements(43), 
          phi_sample_ack => loadKernelChannel_CP_1635_elements(44), 
          phi_update_req => loadKernelChannel_CP_1635_elements(45), 
          phi_update_ack => loadKernelChannel_CP_1635_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_1635_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1773_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_1635_elements(16);
        preds(1)  <= loadKernelChannel_CP_1635_elements(17);
        entry_tmerge_1773 : transition_merge -- 
          generic map(name => " entry_tmerge_1773")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_1635_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_594_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_643_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_607_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_652_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_652_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_652_wire : std_logic_vector(63 downto 0);
    signal NOT_u1_u1_617_wire : std_logic_vector(0 downto 0);
    signal R_sh_start_541_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_541_scaled : std_logic_vector(13 downto 0);
    signal SHL_u16_u16_530_wire : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_559_wire : std_logic_vector(15 downto 0);
    signal SUB_u64_u64_595_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_680_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_620_wire : std_logic_vector(0 downto 0);
    signal ULT_u64_u1_681_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_542_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_542_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_653_root_address : std_logic_vector(13 downto 0);
    signal ea1_554 : std_logic_vector(63 downto 0);
    signal ea2_562 : std_logic_vector(63 downto 0);
    signal ea3_568 : std_logic_vector(63 downto 0);
    signal fetch_addr_544 : std_logic_vector(31 downto 0);
    signal fetch_addr_655 : std_logic_vector(31 downto 0);
    signal fetch_val_585 : std_logic_vector(63 downto 0);
    signal fetch_val_616_delayed_13_0_669 : std_logic_vector(63 downto 0);
    signal first_fill_573 : std_logic_vector(0 downto 0);
    signal fn_608_delayed_7_0_658 : std_logic_vector(0 downto 0);
    signal fn_614_delayed_13_0_666 : std_logic_vector(0 downto 0);
    signal fn_646 : std_logic_vector(0 downto 0);
    signal fv_663 : std_logic_vector(63 downto 0);
    signal konst_529_wire_constant : std_logic_vector(15 downto 0);
    signal konst_535_wire_constant : std_logic_vector(63 downto 0);
    signal konst_558_wire_constant : std_logic_vector(15 downto 0);
    signal konst_571_wire_constant : std_logic_vector(63 downto 0);
    signal konst_591_wire_constant : std_logic_vector(63 downto 0);
    signal konst_593_wire_constant : std_logic_vector(63 downto 0);
    signal konst_596_wire_constant : std_logic_vector(63 downto 0);
    signal konst_601_wire_constant : std_logic_vector(63 downto 0);
    signal konst_642_wire_constant : std_logic_vector(63 downto 0);
    signal konst_644_wire_constant : std_logic_vector(63 downto 0);
    signal konst_651_wire_constant : std_logic_vector(63 downto 0);
    signal konst_679_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_548 : std_logic_vector(63 downto 0);
    signal my_fetch_548_587_buffered : std_logic_vector(63 downto 0);
    signal my_num1_598 : std_logic_vector(63 downto 0);
    signal mycount_581 : std_logic_vector(63 downto 0);
    signal nfetch_val_675 : std_logic_vector(63 downto 0);
    signal nfetch_val_675_588_buffered : std_logic_vector(63 downto 0);
    signal nmycount_603 : std_logic_vector(63 downto 0);
    signal nmycount_603_584_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_547_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_547_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_547_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_547_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_547_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_662_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_662_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_662_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_662_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_662_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_size_532 : std_logic_vector(15 downto 0);
    signal send_to_1_614 : std_logic_vector(0 downto 0);
    signal send_to_2_622 : std_logic_vector(0 downto 0);
    signal send_to_3_627 : std_logic_vector(0 downto 0);
    signal sh_start_537 : std_logic_vector(63 downto 0);
    signal start_add_583_buffered : std_logic_vector(63 downto 0);
    signal start_next_577 : std_logic_vector(7 downto 0);
    signal type_cast_552_wire : std_logic_vector(63 downto 0);
    signal type_cast_560_wire : std_logic_vector(63 downto 0);
    signal type_cast_566_wire : std_logic_vector(63 downto 0);
    signal var_val_609 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_542_constant_part_of_offset <= "00000000000000";
    array_obj_ref_542_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_542_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_542_resized_base_address <= "00000000000000";
    array_obj_ref_653_constant_part_of_offset <= "00000000000000";
    array_obj_ref_653_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_653_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_653_resized_base_address <= "00000000000000";
    konst_529_wire_constant <= "0000000000000001";
    konst_535_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_558_wire_constant <= "0000000000000001";
    konst_571_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_591_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_593_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_596_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_601_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_642_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_644_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_651_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_679_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_547_word_offset_0 <= "00000000000000";
    ptr_deref_662_word_offset_0 <= "00000000000000";
    phi_stmt_581: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= start_add_583_buffered & nmycount_603_584_buffered;
      req <= phi_stmt_581_req_0 & phi_stmt_581_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_581",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_581_ack_0,
          idata => idata,
          odata => mycount_581,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_581
    phi_stmt_585: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= my_fetch_548_587_buffered & nfetch_val_675_588_buffered;
      req <= phi_stmt_585_req_0 & phi_stmt_585_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_585",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_585_ack_0,
          idata => idata,
          odata => fetch_val_585,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_585
    -- flow-through select operator MUX_674_inst
    nfetch_val_675 <= fv_663 when (fn_614_delayed_13_0_666(0) /=  '0') else fetch_val_616_delayed_13_0_669;
    W_fetch_val_616_delayed_13_0_667_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_616_delayed_13_0_667_inst_req_0;
      W_fetch_val_616_delayed_13_0_667_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_616_delayed_13_0_667_inst_req_1;
      W_fetch_val_616_delayed_13_0_667_inst_ack_1<= rack(0);
      W_fetch_val_616_delayed_13_0_667_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_616_delayed_13_0_667_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_585,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_616_delayed_13_0_669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_608_delayed_7_0_656_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_608_delayed_7_0_656_inst_req_0;
      W_fn_608_delayed_7_0_656_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_608_delayed_7_0_656_inst_req_1;
      W_fn_608_delayed_7_0_656_inst_ack_1<= rack(0);
      W_fn_608_delayed_7_0_656_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_608_delayed_7_0_656_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_608_delayed_7_0_658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_614_delayed_13_0_664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_614_delayed_13_0_664_inst_req_0;
      W_fn_614_delayed_13_0_664_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_614_delayed_13_0_664_inst_req_1;
      W_fn_614_delayed_13_0_664_inst_ack_1<= rack(0);
      W_fn_614_delayed_13_0_664_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_614_delayed_13_0_664_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_614_delayed_13_0_666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_543_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_543_final_reg_req_0;
      addr_of_543_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_543_final_reg_req_1;
      addr_of_543_final_reg_ack_1<= rack(0);
      addr_of_543_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_543_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_542_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_654_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_654_final_reg_req_0;
      addr_of_654_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_654_final_reg_req_1;
      addr_of_654_final_reg_ack_1<= rack(0);
      addr_of_654_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_654_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_653_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_655,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_548_587_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_548_587_buf_req_0;
      my_fetch_548_587_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_548_587_buf_req_1;
      my_fetch_548_587_buf_ack_1<= rack(0);
      my_fetch_548_587_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_548_587_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_548_587_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_675_588_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_675_588_buf_req_0;
      nfetch_val_675_588_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_675_588_buf_req_1;
      nfetch_val_675_588_buf_ack_1<= rack(0);
      nfetch_val_675_588_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_675_588_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_675,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_675_588_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_603_584_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_603_584_buf_req_0;
      nmycount_603_584_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_603_584_buf_req_1;
      nmycount_603_584_buf_ack_1<= rack(0);
      nmycount_603_584_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_603_584_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_603,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_603_584_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_583_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_583_buf_req_0;
      start_add_583_buf_ack_0<= wack(0);
      rreq(0) <= start_add_583_buf_req_1;
      start_add_583_buf_ack_1<= rack(0);
      start_add_583_buf : InterlockBuffer generic map ( -- 
        name => "start_add_583_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_583_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_552_inst
    process(row_size_532) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_532(15 downto 0);
      type_cast_552_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_560_inst
    process(SHL_u16_u16_559_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := SHL_u16_u16_559_wire(15 downto 0);
      type_cast_560_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_566_inst
    process(row_size_532) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_532(15 downto 0);
      type_cast_566_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_608_inst
    process(LSHR_u64_u64_607_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_607_wire(15 downto 0);
      var_val_609 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_542_index_1_rename
    process(R_sh_start_541_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_541_resized;
      ov(13 downto 0) := iv;
      R_sh_start_541_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_542_index_1_resize
    process(sh_start_537) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_537;
      ov := iv(13 downto 0);
      R_sh_start_541_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_542_root_address_inst
    process(array_obj_ref_542_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_542_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_542_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_index_1_rename
    process(LSHR_u64_u64_652_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_652_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_652_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_index_1_resize
    process(LSHR_u64_u64_652_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_652_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_652_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_653_root_address_inst
    process(array_obj_ref_653_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_653_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_653_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_547_addr_0
    process(ptr_deref_547_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_547_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_547_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_547_base_resize
    process(fetch_addr_544) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_544;
      ov := iv(13 downto 0);
      ptr_deref_547_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_547_gather_scatter
    process(ptr_deref_547_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_547_data_0;
      ov(63 downto 0) := iv;
      my_fetch_548 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_547_root_address_inst
    process(ptr_deref_547_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_547_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_547_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_662_addr_0
    process(ptr_deref_662_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_662_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_662_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_662_base_resize
    process(fetch_addr_655) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_655;
      ov := iv(13 downto 0);
      ptr_deref_662_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_662_gather_scatter
    process(ptr_deref_662_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_662_data_0;
      ov(63 downto 0) := iv;
      fv_663 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_662_root_address_inst
    process(ptr_deref_662_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_662_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_662_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_579_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_681_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_579_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_579_branch_req_0,
          ack0 => do_while_stmt_579_branch_ack_0,
          ack1 => do_while_stmt_579_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_531_inst
    process(num_chl_buffer, SHL_u16_u16_530_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_chl_buffer, SHL_u16_u16_530_wire, tmp_var);
      row_size_532 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_553_inst
    process(start_add_buffer, type_cast_552_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_552_wire, tmp_var);
      ea1_554 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_561_inst
    process(start_add_buffer, type_cast_560_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_560_wire, tmp_var);
      ea2_562 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_567_inst
    process(ea2_562, type_cast_566_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ea2_562, type_cast_566_wire, tmp_var);
      ea3_568 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_602_inst
    process(mycount_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_581, konst_601_wire_constant, tmp_var);
      nmycount_603 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_621_inst
    process(NOT_u1_u1_617_wire, ULT_u64_u1_620_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_617_wire, ULT_u64_u1_620_wire, tmp_var);
      send_to_2_622 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_594_inst
    process(mycount_581) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_581, konst_593_wire_constant, tmp_var);
      AND_u64_u64_594_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_643_inst
    process(nmycount_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_603, konst_642_wire_constant, tmp_var);
      AND_u64_u64_643_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_572_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_571_wire_constant, tmp_var);
      first_fill_573 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_645_inst
    process(AND_u64_u64_643_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_643_wire, konst_644_wire_constant, tmp_var);
      fn_646 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_536_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_535_wire_constant, tmp_var);
      sh_start_537 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_607_inst
    process(fetch_val_585, my_num1_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_585, my_num1_598, tmp_var);
      LSHR_u64_u64_607_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_652_inst
    process(nmycount_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_603, konst_651_wire_constant, tmp_var);
      LSHR_u64_u64_652_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_617_inst
    process(send_to_1_614) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", send_to_1_614, tmp_var);
      NOT_u1_u1_617_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u16_u16_530_inst
    process(num_chl_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(num_chl_buffer, konst_529_wire_constant, tmp_var);
      SHL_u16_u16_530_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_559_inst
    process(row_size_532) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(row_size_532, konst_558_wire_constant, tmp_var);
      SHL_u16_u16_559_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_597_inst
    process(SUB_u64_u64_595_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_595_wire, konst_596_wire_constant, tmp_var);
      my_num1_598 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_595_inst
    process(konst_591_wire_constant, AND_u64_u64_594_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_591_wire_constant, AND_u64_u64_594_wire, tmp_var);
      SUB_u64_u64_595_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_680_inst
    process(ea3_568) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(ea3_568, konst_679_wire_constant, tmp_var);
      SUB_u64_u64_680_wire <= tmp_var; --
    end process;
    -- binary operator UGE_u64_u1_626_inst
    process(mycount_581, ea2_562) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(mycount_581, ea2_562, tmp_var);
      send_to_3_627 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_613_inst
    process(mycount_581, ea1_554) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_581, ea1_554, tmp_var);
      send_to_1_614 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_620_inst
    process(mycount_581, ea2_562) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_581, ea2_562, tmp_var);
      ULT_u64_u1_620_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_681_inst
    process(mycount_581, SUB_u64_u64_680_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_581, SUB_u64_u64_680_wire, tmp_var);
      ULT_u64_u1_681_wire <= tmp_var; --
    end process;
    -- shared split operator group (23) : array_obj_ref_542_index_offset 
    ApIntAdd_group_23: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_541_scaled;
      array_obj_ref_542_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_542_index_offset_req_0;
      array_obj_ref_542_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_542_index_offset_req_1;
      array_obj_ref_542_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_23_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : array_obj_ref_653_index_offset 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_652_scaled;
      array_obj_ref_653_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_653_index_offset_req_0;
      array_obj_ref_653_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_653_index_offset_req_1;
      array_obj_ref_653_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared load operator group (0) : ptr_deref_547_load_0 ptr_deref_662_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_547_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_662_load_0_req_0;
      ptr_deref_547_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_662_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_547_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_662_load_0_req_1;
      ptr_deref_547_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_662_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_608_delayed_7_0_658(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_547_word_address_0 & ptr_deref_662_word_address_0;
      ptr_deref_547_data_0 <= data_out(127 downto 64);
      ptr_deref_662_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_576_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_576_inst_req_0;
      RPIPE_input_done_pipe_576_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_576_inst_req_1;
      RPIPE_input_done_pipe_576_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_573(0);
      start_next_577 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_629_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_629_inst_req_0;
      WPIPE_kernel_pipe1_629_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_629_inst_req_1;
      WPIPE_kernel_pipe1_629_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_614(0);
      data_in <= var_val_609;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe2_633_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_633_inst_req_0;
      WPIPE_kernel_pipe2_633_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_633_inst_req_1;
      WPIPE_kernel_pipe2_633_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_622(0);
      data_in <= var_val_609;
      kernel_pipe2_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_kernel_pipe3_637_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe3_637_inst_req_0;
      WPIPE_kernel_pipe3_637_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe3_637_inst_req_1;
      WPIPE_kernel_pipe3_637_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_627(0);
      data_in <= var_val_609;
      kernel_pipe3_write_2_gI: SplitGuardInterface generic map(name => "kernel_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "kernel_pipe3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe3_pipe_write_req(0),
          oack => kernel_pipe3_pipe_write_ack(0),
          odata => kernel_pipe3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_size_pipe_683_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_683_inst_req_0;
      WPIPE_size_pipe_683_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_683_inst_req_1;
      WPIPE_size_pipe_683_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= num_chl_buffer;
      size_pipe_write_3_gI: SplitGuardInterface generic map(name => "size_pipe_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_3: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(63 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_2093_start: Boolean;
  signal sendB_CP_2093_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_702_branch_ack_0 : boolean;
  signal ptr_deref_998_store_0_ack_0 : boolean;
  signal if_stmt_702_branch_ack_1 : boolean;
  signal array_obj_ref_748_index_offset_req_1 : boolean;
  signal array_obj_ref_748_index_offset_ack_1 : boolean;
  signal array_obj_ref_748_index_offset_req_0 : boolean;
  signal type_cast_1009_inst_ack_0 : boolean;
  signal type_cast_1051_inst_ack_0 : boolean;
  signal array_obj_ref_1140_final_reg_ack_0 : boolean;
  signal type_cast_1009_inst_req_1 : boolean;
  signal if_stmt_702_branch_req_0 : boolean;
  signal array_obj_ref_748_index_offset_ack_0 : boolean;
  signal array_obj_ref_1128_final_reg_req_0 : boolean;
  signal array_obj_ref_1128_final_reg_ack_0 : boolean;
  signal type_cast_1009_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1146_inst_ack_1 : boolean;
  signal array_obj_ref_1140_final_reg_req_1 : boolean;
  signal type_cast_1051_inst_req_1 : boolean;
  signal array_obj_ref_1128_index_offset_req_0 : boolean;
  signal ptr_deref_1061_store_0_req_0 : boolean;
  signal array_obj_ref_1128_index_offset_ack_0 : boolean;
  signal ptr_deref_1061_store_0_ack_0 : boolean;
  signal array_obj_ref_1140_final_reg_ack_1 : boolean;
  signal type_cast_1051_inst_ack_1 : boolean;
  signal ptr_deref_1019_store_0_req_0 : boolean;
  signal ptr_deref_1151_load_0_req_1 : boolean;
  signal ptr_deref_1151_load_0_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1146_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1146_inst_ack_0 : boolean;
  signal ptr_deref_1040_store_0_req_0 : boolean;
  signal ptr_deref_1019_store_0_ack_0 : boolean;
  signal ptr_deref_1144_load_0_req_1 : boolean;
  signal array_obj_ref_1128_index_offset_req_1 : boolean;
  signal array_obj_ref_1140_index_offset_req_0 : boolean;
  signal array_obj_ref_1140_index_offset_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1146_inst_req_1 : boolean;
  signal ptr_deref_1144_load_0_req_0 : boolean;
  signal ptr_deref_1144_load_0_ack_1 : boolean;
  signal ptr_deref_998_store_0_req_1 : boolean;
  signal ptr_deref_1040_store_0_ack_0 : boolean;
  signal addr_of_749_final_reg_req_0 : boolean;
  signal addr_of_749_final_reg_ack_0 : boolean;
  signal addr_of_749_final_reg_req_1 : boolean;
  signal addr_of_749_final_reg_ack_1 : boolean;
  signal ptr_deref_753_load_0_req_0 : boolean;
  signal ptr_deref_753_load_0_ack_0 : boolean;
  signal ptr_deref_753_load_0_req_1 : boolean;
  signal ptr_deref_753_load_0_ack_1 : boolean;
  signal type_cast_757_inst_req_0 : boolean;
  signal type_cast_757_inst_ack_0 : boolean;
  signal type_cast_757_inst_req_1 : boolean;
  signal type_cast_757_inst_ack_1 : boolean;
  signal type_cast_767_inst_req_0 : boolean;
  signal type_cast_767_inst_ack_0 : boolean;
  signal type_cast_767_inst_req_1 : boolean;
  signal type_cast_767_inst_ack_1 : boolean;
  signal type_cast_777_inst_req_0 : boolean;
  signal type_cast_777_inst_ack_0 : boolean;
  signal type_cast_777_inst_req_1 : boolean;
  signal type_cast_777_inst_ack_1 : boolean;
  signal type_cast_787_inst_req_0 : boolean;
  signal type_cast_787_inst_ack_0 : boolean;
  signal type_cast_787_inst_req_1 : boolean;
  signal type_cast_787_inst_ack_1 : boolean;
  signal type_cast_797_inst_req_0 : boolean;
  signal type_cast_797_inst_ack_0 : boolean;
  signal type_cast_797_inst_req_1 : boolean;
  signal type_cast_797_inst_ack_1 : boolean;
  signal type_cast_807_inst_req_0 : boolean;
  signal type_cast_807_inst_ack_0 : boolean;
  signal type_cast_807_inst_req_1 : boolean;
  signal type_cast_807_inst_ack_1 : boolean;
  signal type_cast_817_inst_req_0 : boolean;
  signal type_cast_817_inst_ack_0 : boolean;
  signal type_cast_817_inst_req_1 : boolean;
  signal type_cast_817_inst_ack_1 : boolean;
  signal type_cast_827_inst_req_0 : boolean;
  signal type_cast_827_inst_ack_0 : boolean;
  signal type_cast_827_inst_req_1 : boolean;
  signal type_cast_827_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_829_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_829_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_829_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_829_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_832_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_832_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_832_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_832_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_835_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_835_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_835_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_835_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_838_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_838_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_838_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_838_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_841_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_841_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_841_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_841_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_844_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_844_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_844_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_844_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_847_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_847_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_847_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_847_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_850_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_850_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_850_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_850_inst_ack_1 : boolean;
  signal type_cast_1051_inst_req_0 : boolean;
  signal if_stmt_864_branch_req_0 : boolean;
  signal array_obj_ref_1140_final_reg_req_0 : boolean;
  signal ptr_deref_998_store_0_req_0 : boolean;
  signal if_stmt_864_branch_ack_1 : boolean;
  signal if_stmt_864_branch_ack_0 : boolean;
  signal type_cast_1009_inst_req_0 : boolean;
  signal if_stmt_916_branch_req_0 : boolean;
  signal if_stmt_916_branch_ack_1 : boolean;
  signal if_stmt_916_branch_ack_0 : boolean;
  signal type_cast_925_inst_req_0 : boolean;
  signal type_cast_925_inst_ack_0 : boolean;
  signal type_cast_925_inst_req_1 : boolean;
  signal type_cast_925_inst_ack_1 : boolean;
  signal ptr_deref_1151_load_0_ack_0 : boolean;
  signal if_stmt_1070_branch_ack_0 : boolean;
  signal ptr_deref_1040_store_0_ack_1 : boolean;
  signal ptr_deref_1040_store_0_req_1 : boolean;
  signal array_obj_ref_931_index_offset_req_0 : boolean;
  signal array_obj_ref_931_index_offset_ack_0 : boolean;
  signal array_obj_ref_931_index_offset_req_1 : boolean;
  signal array_obj_ref_931_index_offset_ack_1 : boolean;
  signal ptr_deref_1144_load_0_ack_0 : boolean;
  signal array_obj_ref_1140_index_offset_ack_1 : boolean;
  signal addr_of_932_final_reg_req_0 : boolean;
  signal addr_of_932_final_reg_ack_0 : boolean;
  signal addr_of_932_final_reg_req_1 : boolean;
  signal addr_of_932_final_reg_ack_1 : boolean;
  signal ptr_deref_1151_load_0_req_0 : boolean;
  signal if_stmt_1070_branch_ack_1 : boolean;
  signal if_stmt_1070_branch_req_0 : boolean;
  signal ptr_deref_936_load_0_req_0 : boolean;
  signal type_cast_1030_inst_ack_1 : boolean;
  signal ptr_deref_936_load_0_ack_0 : boolean;
  signal ptr_deref_936_load_0_req_1 : boolean;
  signal type_cast_1030_inst_req_1 : boolean;
  signal ptr_deref_936_load_0_ack_1 : boolean;
  signal type_cast_946_inst_req_0 : boolean;
  signal type_cast_946_inst_ack_0 : boolean;
  signal array_obj_ref_1128_final_reg_ack_1 : boolean;
  signal type_cast_946_inst_req_1 : boolean;
  signal type_cast_946_inst_ack_1 : boolean;
  signal array_obj_ref_1128_index_offset_ack_1 : boolean;
  signal ptr_deref_1061_store_0_ack_1 : boolean;
  signal ptr_deref_1061_store_0_req_1 : boolean;
  signal type_cast_1030_inst_ack_0 : boolean;
  signal type_cast_1030_inst_req_0 : boolean;
  signal array_obj_ref_1128_final_reg_req_1 : boolean;
  signal ptr_deref_956_store_0_req_0 : boolean;
  signal ptr_deref_956_store_0_ack_0 : boolean;
  signal ptr_deref_956_store_0_req_1 : boolean;
  signal ptr_deref_956_store_0_ack_1 : boolean;
  signal array_obj_ref_1140_index_offset_req_1 : boolean;
  signal ptr_deref_1019_store_0_ack_1 : boolean;
  signal ptr_deref_1019_store_0_req_1 : boolean;
  signal type_cast_967_inst_req_0 : boolean;
  signal type_cast_967_inst_ack_0 : boolean;
  signal type_cast_967_inst_req_1 : boolean;
  signal type_cast_967_inst_ack_1 : boolean;
  signal ptr_deref_998_store_0_ack_1 : boolean;
  signal ptr_deref_977_store_0_req_0 : boolean;
  signal ptr_deref_977_store_0_ack_0 : boolean;
  signal ptr_deref_977_store_0_req_1 : boolean;
  signal ptr_deref_977_store_0_ack_1 : boolean;
  signal type_cast_988_inst_req_0 : boolean;
  signal type_cast_988_inst_ack_0 : boolean;
  signal type_cast_988_inst_req_1 : boolean;
  signal type_cast_988_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1153_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1153_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1153_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1153_inst_ack_1 : boolean;
  signal if_stmt_1167_branch_req_0 : boolean;
  signal if_stmt_1167_branch_ack_1 : boolean;
  signal if_stmt_1167_branch_ack_0 : boolean;
  signal phi_stmt_736_req_0 : boolean;
  signal type_cast_742_inst_req_0 : boolean;
  signal type_cast_742_inst_ack_0 : boolean;
  signal type_cast_742_inst_req_1 : boolean;
  signal type_cast_742_inst_ack_1 : boolean;
  signal phi_stmt_736_req_1 : boolean;
  signal phi_stmt_736_ack_0 : boolean;
  signal phi_stmt_896_req_1 : boolean;
  signal type_cast_899_inst_req_0 : boolean;
  signal type_cast_899_inst_ack_0 : boolean;
  signal type_cast_899_inst_req_1 : boolean;
  signal type_cast_899_inst_ack_1 : boolean;
  signal phi_stmt_896_req_0 : boolean;
  signal phi_stmt_896_ack_0 : boolean;
  signal phi_stmt_1110_req_0 : boolean;
  signal type_cast_1116_inst_req_0 : boolean;
  signal type_cast_1116_inst_ack_0 : boolean;
  signal type_cast_1116_inst_req_1 : boolean;
  signal type_cast_1116_inst_ack_1 : boolean;
  signal phi_stmt_1110_req_1 : boolean;
  signal phi_stmt_1110_ack_0 : boolean;
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(2 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= size;
  size_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_2093_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2093_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_2093_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2093_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_2093: Block -- control-path 
    signal sendB_CP_2093_elements: BooleanArray(137 downto 0);
    -- 
  begin -- 
    sendB_CP_2093_elements(0) <= sendB_CP_2093_start;
    sendB_CP_2093_symbol <= sendB_CP_2093_elements(137);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_else_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/assign_stmt_695_to_assign_stmt_701/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/assign_stmt_695_to_assign_stmt_701/$exit
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/R_cmp77_703_place
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_689/$entry
      -- CP-element group 0: 	 branch_block_stmt_689/branch_block_stmt_689__entry__
      -- CP-element group 0: 	 branch_block_stmt_689/assign_stmt_695_to_assign_stmt_701__entry__
      -- CP-element group 0: 	 branch_block_stmt_689/assign_stmt_695_to_assign_stmt_701__exit__
      -- CP-element group 0: 	 branch_block_stmt_689/if_stmt_702__entry__
      -- 
    branch_req_2157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(0), ack => if_stmt_702_branch_req_0); -- 
    -- CP-element group 1:  merge  transition  place  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	119 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_689/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_733/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/if_stmt_702_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_689/if_stmt_702_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_689/bbx_xnph_forx_xbody
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_733/$exit
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708__exit__
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_733__entry__
      -- CP-element group 1: 	 branch_block_stmt_689/assign_stmt_714_to_assign_stmt_733__exit__
      -- CP-element group 1: 	 branch_block_stmt_689/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_689/merge_stmt_708_PhiAck/dummy
      -- CP-element group 1: 	 branch_block_stmt_689/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/bbx_xnph_forx_xbody_PhiReq/phi_stmt_736/$entry
      -- CP-element group 1: 	 branch_block_stmt_689/bbx_xnph_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/$entry
      -- 
    if_choice_transition_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_702_branch_ack_1, ack => sendB_CP_2093_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	125 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_689/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_689/if_stmt_702_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_689/if_stmt_702_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_896/$entry
      -- CP-element group 2: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/$entry
      -- 
    else_choice_transition_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_702_branch_ack_0, ack => sendB_CP_2093_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	124 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	48 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_sample_complete
      -- CP-element group 3: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_Sample/$exit
      -- 
    ack_2200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_748_index_offset_ack_0, ack => sendB_CP_2093_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	124 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (11) 
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_offset_calculated
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_Update/ack
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_root_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_base_plus_offset/$entry
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_base_plus_offset/$exit
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_request/$entry
      -- CP-element group 4: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_request/req
      -- 
    ack_2205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_748_index_offset_ack_1, ack => sendB_CP_2093_elements(4)); -- 
    req_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(4), ack => addr_of_749_final_reg_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_request/$exit
      -- CP-element group 5: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_request/ack
      -- 
    ack_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_749_final_reg_ack_0, ack => sendB_CP_2093_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	124 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (24) 
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_complete/ack
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_word_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_address_resized
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_addr_resize/$entry
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_addr_resize/$exit
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_addr_resize/base_resize_req
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_addr_resize/base_resize_ack
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_word_addrgen/$entry
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_word_addrgen/$exit
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_word_addrgen/root_register_req
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_word_addrgen/root_register_ack
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Sample/word_access_start/$entry
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Sample/word_access_start/word_0/$entry
      -- CP-element group 6: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Sample/word_access_start/word_0/rr
      -- 
    ack_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_749_final_reg_ack_1, ack => sendB_CP_2093_elements(6)); -- 
    rr_2253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(6), ack => ptr_deref_753_load_0_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Sample/word_access_start/word_0/ra
      -- 
    ra_2254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_753_load_0_ack_0, ack => sendB_CP_2093_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	124 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	11 
    -- CP-element group 8: 	13 
    -- CP-element group 8: 	15 
    -- CP-element group 8: 	17 
    -- CP-element group 8: 	19 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (33) 
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/ptr_deref_753_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/ptr_deref_753_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/ptr_deref_753_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/ptr_deref_753_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_Sample/rr
      -- 
    ca_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_753_load_0_ack_1, ack => sendB_CP_2093_elements(8)); -- 
    rr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => type_cast_757_inst_req_0); -- 
    rr_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => type_cast_767_inst_req_0); -- 
    rr_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => type_cast_777_inst_req_0); -- 
    rr_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => type_cast_787_inst_req_0); -- 
    rr_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => type_cast_797_inst_req_0); -- 
    rr_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => type_cast_807_inst_req_0); -- 
    rr_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => type_cast_817_inst_req_0); -- 
    rr_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(8), ack => type_cast_827_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_Sample/ra
      -- 
    ra_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_757_inst_ack_0, ack => sendB_CP_2093_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	124 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	45 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_Update/ca
      -- 
    ca_2284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_757_inst_ack_1, ack => sendB_CP_2093_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_Sample/ra
      -- 
    ra_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_767_inst_ack_0, ack => sendB_CP_2093_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	124 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	42 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_Update/ca
      -- 
    ca_2298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_767_inst_ack_1, ack => sendB_CP_2093_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_Sample/ra
      -- 
    ra_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_777_inst_ack_0, ack => sendB_CP_2093_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	124 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	39 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_Update/ca
      -- 
    ca_2312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_777_inst_ack_1, ack => sendB_CP_2093_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	8 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_Sample/ra
      -- 
    ra_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_787_inst_ack_0, ack => sendB_CP_2093_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	124 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	36 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_Update/ca
      -- 
    ca_2326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_787_inst_ack_1, ack => sendB_CP_2093_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	8 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_Sample/ra
      -- 
    ra_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_0, ack => sendB_CP_2093_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	124 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_Update/ca
      -- 
    ca_2340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_1, ack => sendB_CP_2093_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	8 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_Sample/ra
      -- 
    ra_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_0, ack => sendB_CP_2093_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	124 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	30 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_Update/ca
      -- 
    ca_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_1, ack => sendB_CP_2093_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_Sample/ra
      -- 
    ra_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_0, ack => sendB_CP_2093_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	124 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_Update/ca
      -- 
    ca_2368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_1, ack => sendB_CP_2093_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_Sample/ra
      -- 
    ra_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_0, ack => sendB_CP_2093_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	124 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_Sample/req
      -- 
    ca_2382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_827_inst_ack_1, ack => sendB_CP_2093_elements(24)); -- 
    req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(24), ack => WPIPE_maxpool_output_pipe_829_inst_req_0); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_update_start_
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_Sample/ack
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_Update/req
      -- 
    ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_829_inst_ack_0, ack => sendB_CP_2093_elements(25)); -- 
    req_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(25), ack => WPIPE_maxpool_output_pipe_829_inst_req_1); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_829_Update/ack
      -- 
    ack_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_829_inst_ack_1, ack => sendB_CP_2093_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: 	22 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_Sample/req
      -- 
    req_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(27), ack => WPIPE_maxpool_output_pipe_832_inst_req_0); -- 
    sendB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(26) & sendB_CP_2093_elements(22);
      gj_sendB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_update_start_
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_Update/req
      -- 
    ack_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_832_inst_ack_0, ack => sendB_CP_2093_elements(28)); -- 
    req_2409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(28), ack => WPIPE_maxpool_output_pipe_832_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_832_Update/ack
      -- 
    ack_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_832_inst_ack_1, ack => sendB_CP_2093_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: 	20 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_Sample/req
      -- 
    req_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(30), ack => WPIPE_maxpool_output_pipe_835_inst_req_0); -- 
    sendB_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(29) & sendB_CP_2093_elements(20);
      gj_sendB_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_update_start_
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_Update/req
      -- 
    ack_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_835_inst_ack_0, ack => sendB_CP_2093_elements(31)); -- 
    req_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(31), ack => WPIPE_maxpool_output_pipe_835_inst_req_1); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_835_Update/ack
      -- 
    ack_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_835_inst_ack_1, ack => sendB_CP_2093_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	18 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_Sample/req
      -- 
    req_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(33), ack => WPIPE_maxpool_output_pipe_838_inst_req_0); -- 
    sendB_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(32) & sendB_CP_2093_elements(18);
      gj_sendB_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_update_start_
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_Update/req
      -- 
    ack_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_838_inst_ack_0, ack => sendB_CP_2093_elements(34)); -- 
    req_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(34), ack => WPIPE_maxpool_output_pipe_838_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_838_Update/ack
      -- 
    ack_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_838_inst_ack_1, ack => sendB_CP_2093_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	16 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_Sample/req
      -- 
    req_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(36), ack => WPIPE_maxpool_output_pipe_841_inst_req_0); -- 
    sendB_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(35) & sendB_CP_2093_elements(16);
      gj_sendB_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_update_start_
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_Update/req
      -- 
    ack_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_841_inst_ack_0, ack => sendB_CP_2093_elements(37)); -- 
    req_2451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(37), ack => WPIPE_maxpool_output_pipe_841_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_841_Update/ack
      -- 
    ack_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_841_inst_ack_1, ack => sendB_CP_2093_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: 	14 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_Sample/req
      -- 
    req_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(39), ack => WPIPE_maxpool_output_pipe_844_inst_req_0); -- 
    sendB_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(38) & sendB_CP_2093_elements(14);
      gj_sendB_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_update_start_
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_Update/req
      -- 
    ack_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_844_inst_ack_0, ack => sendB_CP_2093_elements(40)); -- 
    req_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(40), ack => WPIPE_maxpool_output_pipe_844_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_844_Update/ack
      -- 
    ack_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_844_inst_ack_1, ack => sendB_CP_2093_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	12 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_Sample/req
      -- 
    req_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(42), ack => WPIPE_maxpool_output_pipe_847_inst_req_0); -- 
    sendB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(41) & sendB_CP_2093_elements(12);
      gj_sendB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_update_start_
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_Update/req
      -- 
    ack_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_847_inst_ack_0, ack => sendB_CP_2093_elements(43)); -- 
    req_2479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(43), ack => WPIPE_maxpool_output_pipe_847_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_847_Update/ack
      -- 
    ack_2480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_847_inst_ack_1, ack => sendB_CP_2093_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_Sample/req
      -- 
    req_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(45), ack => WPIPE_maxpool_output_pipe_850_inst_req_0); -- 
    sendB_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(44) & sendB_CP_2093_elements(10);
      gj_sendB_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_update_start_
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_Update/req
      -- 
    ack_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_850_inst_ack_0, ack => sendB_CP_2093_elements(46)); -- 
    req_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(46), ack => WPIPE_maxpool_output_pipe_850_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/WPIPE_maxpool_output_pipe_850_Update/ack
      -- 
    ack_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_850_inst_ack_1, ack => sendB_CP_2093_elements(47)); -- 
    -- CP-element group 48:  branch  join  transition  place  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	3 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (10) 
      -- CP-element group 48: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863__exit__
      -- CP-element group 48: 	 branch_block_stmt_689/if_stmt_864__entry__
      -- CP-element group 48: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/$exit
      -- CP-element group 48: 	 branch_block_stmt_689/if_stmt_864_dead_link/$entry
      -- CP-element group 48: 	 branch_block_stmt_689/if_stmt_864_eval_test/$entry
      -- CP-element group 48: 	 branch_block_stmt_689/if_stmt_864_eval_test/$exit
      -- CP-element group 48: 	 branch_block_stmt_689/if_stmt_864_eval_test/branch_req
      -- CP-element group 48: 	 branch_block_stmt_689/R_exitcond_865_place
      -- CP-element group 48: 	 branch_block_stmt_689/if_stmt_864_if_link/$entry
      -- CP-element group 48: 	 branch_block_stmt_689/if_stmt_864_else_link/$entry
      -- 
    branch_req_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(48), ack => if_stmt_864_branch_req_0); -- 
    sendB_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(47) & sendB_CP_2093_elements(3);
      gj_sendB_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	126 
    -- CP-element group 49: 	127 
    -- CP-element group 49:  members (24) 
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 49: 	 branch_block_stmt_689/assign_stmt_877_to_assign_stmt_893__exit__
      -- CP-element group 49: 	 branch_block_stmt_689/assign_stmt_877_to_assign_stmt_893__entry__
      -- CP-element group 49: 	 branch_block_stmt_689/merge_stmt_870__exit__
      -- CP-element group 49: 	 branch_block_stmt_689/if_stmt_864_if_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_689/if_stmt_864_if_link/if_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 49: 	 branch_block_stmt_689/assign_stmt_877_to_assign_stmt_893/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/assign_stmt_877_to_assign_stmt_893/$exit
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 49: 	 branch_block_stmt_689/merge_stmt_870_PhiReqMerge
      -- CP-element group 49: 	 branch_block_stmt_689/merge_stmt_870_PhiAck/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/merge_stmt_870_PhiAck/$exit
      -- CP-element group 49: 	 branch_block_stmt_689/merge_stmt_870_PhiAck/dummy
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_864_branch_ack_1, ack => sendB_CP_2093_elements(49)); -- 
    rr_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(49), ack => type_cast_899_inst_req_0); -- 
    cr_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(49), ack => type_cast_899_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  place  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	120 
    -- CP-element group 50: 	121 
    -- CP-element group 50:  members (12) 
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_864_else_link/$exit
      -- CP-element group 50: 	 branch_block_stmt_689/if_stmt_864_else_link/else_choice_transition
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_864_branch_ack_0, ack => sendB_CP_2093_elements(50)); -- 
    rr_3348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(50), ack => type_cast_742_inst_req_0); -- 
    cr_3353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(50), ack => type_cast_742_inst_req_1); -- 
    -- CP-element group 51:  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	130 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	137 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_689/if_stmt_916_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_689/if_stmt_916_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_689/forx_xend_sendRemainingElementsx_xexit
      -- CP-element group 51: 	 branch_block_stmt_689/forx_xend_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_689/forx_xend_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_916_branch_ack_1, ack => sendB_CP_2093_elements(51)); -- 
    -- CP-element group 52:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	130 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	70 
    -- CP-element group 52: 	65 
    -- CP-element group 52: 	72 
    -- CP-element group 52: 	67 
    -- CP-element group 52: 	68 
    -- CP-element group 52: 	73 
    -- CP-element group 52: 	75 
    -- CP-element group 52: 	77 
    -- CP-element group 52: 	78 
    -- CP-element group 52: 	80 
    -- CP-element group 52: 	82 
    -- CP-element group 52: 	83 
    -- CP-element group 52: 	85 
    -- CP-element group 52: 	87 
    -- CP-element group 52: 	88 
    -- CP-element group 52: 	90 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52: 	56 
    -- CP-element group 52: 	58 
    -- CP-element group 52: 	60 
    -- CP-element group 52: 	62 
    -- CP-element group 52: 	63 
    -- CP-element group 52:  members (186) 
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069__entry__
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/merge_stmt_922__exit__
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/if_stmt_916_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/if_stmt_916_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xend_ifx_xthen
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_resized_1
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_scaled_1
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_computed_1
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_resize_1/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_resize_1/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_resize_1/index_resize_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_resize_1/index_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_scale_1/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_scale_1/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_scale_1/scale_rename_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_index_scale_1/scale_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_update_start
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_Update/req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_complete/req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Update/word_access_complete/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Update/word_access_complete/word_0/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Update/word_access_complete/word_0/cr
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_update_start_
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_Update/cr
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xend_ifx_xthen_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/forx_xend_ifx_xthen_PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/merge_stmt_922_PhiReqMerge
      -- CP-element group 52: 	 branch_block_stmt_689/merge_stmt_922_PhiAck/$entry
      -- CP-element group 52: 	 branch_block_stmt_689/merge_stmt_922_PhiAck/$exit
      -- CP-element group 52: 	 branch_block_stmt_689/merge_stmt_922_PhiAck/dummy
      -- 
    else_choice_transition_2536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_916_branch_ack_0, ack => sendB_CP_2093_elements(52)); -- 
    cr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_1009_inst_req_1); -- 
    cr_2984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_1051_inst_req_1); -- 
    cr_2842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => ptr_deref_998_store_0_req_1); -- 
    rr_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_925_inst_req_0); -- 
    cr_2554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_925_inst_req_1); -- 
    cr_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => ptr_deref_1040_store_0_req_1); -- 
    req_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => array_obj_ref_931_index_offset_req_0); -- 
    req_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => array_obj_ref_931_index_offset_req_1); -- 
    req_2600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => addr_of_932_final_reg_req_1); -- 
    cr_2645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => ptr_deref_936_load_0_req_1); -- 
    cr_2920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_1030_inst_req_1); -- 
    cr_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_946_inst_req_1); -- 
    cr_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => ptr_deref_1061_store_0_req_1); -- 
    cr_2714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => ptr_deref_956_store_0_req_1); -- 
    cr_2906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => ptr_deref_1019_store_0_req_1); -- 
    cr_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_967_inst_req_1); -- 
    cr_2778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => ptr_deref_977_store_0_req_1); -- 
    cr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(52), ack => type_cast_988_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_Sample/ra
      -- 
    ra_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_925_inst_ack_0, ack => sendB_CP_2093_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	96 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_925_Update/ca
      -- 
    ca_2555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_925_inst_ack_1, ack => sendB_CP_2093_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	96 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_sample_complete
      -- CP-element group 55: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_Sample/ack
      -- 
    ack_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_931_index_offset_ack_0, ack => sendB_CP_2093_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	52 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (11) 
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_offset_calculated
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_final_index_sum_regn_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/array_obj_ref_931_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_request/$entry
      -- CP-element group 56: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_request/req
      -- 
    ack_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_931_index_offset_ack_1, ack => sendB_CP_2093_elements(56)); -- 
    req_2595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(56), ack => addr_of_932_final_reg_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_request/$exit
      -- CP-element group 57: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_request/ack
      -- 
    ack_2596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_932_final_reg_ack_0, ack => sendB_CP_2093_elements(57)); -- 
    -- CP-element group 58:  join  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	52 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_complete/$exit
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/addr_of_932_complete/ack
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_word_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_address_resized
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_addr_resize/$entry
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_addr_resize/$exit
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_addr_resize/base_resize_req
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_addr_resize/base_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_word_addrgen/$entry
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_word_addrgen/$exit
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_word_addrgen/root_register_req
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_word_addrgen/root_register_ack
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Sample/word_access_start/$entry
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Sample/word_access_start/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Sample/word_access_start/word_0/rr
      -- 
    ack_2601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_932_final_reg_ack_1, ack => sendB_CP_2093_elements(58)); -- 
    rr_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(58), ack => ptr_deref_936_load_0_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Sample/word_access_start/$exit
      -- CP-element group 59: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Sample/word_access_start/word_0/$exit
      -- CP-element group 59: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Sample/word_access_start/word_0/ra
      -- 
    ra_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_936_load_0_ack_0, ack => sendB_CP_2093_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	52 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	71 
    -- CP-element group 60: 	66 
    -- CP-element group 60: 	76 
    -- CP-element group 60: 	81 
    -- CP-element group 60: 	86 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (27) 
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/word_access_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/word_access_complete/word_0/$exit
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/word_access_complete/word_0/ca
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/ptr_deref_936_Merge/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/ptr_deref_936_Merge/$exit
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/ptr_deref_936_Merge/merge_req
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_936_Update/ptr_deref_936_Merge/merge_ack
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_Sample/rr
      -- 
    ca_2646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_936_load_0_ack_1, ack => sendB_CP_2093_elements(60)); -- 
    rr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(60), ack => type_cast_988_inst_req_0); -- 
    rr_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(60), ack => type_cast_967_inst_req_0); -- 
    rr_2851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(60), ack => type_cast_1009_inst_req_0); -- 
    rr_2915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(60), ack => type_cast_1030_inst_req_0); -- 
    rr_2979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(60), ack => type_cast_1051_inst_req_0); -- 
    rr_2659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(60), ack => type_cast_946_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_Sample/ra
      -- 
    ra_2660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_946_inst_ack_0, ack => sendB_CP_2093_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	52 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_946_Update/ca
      -- 
    ca_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_946_inst_ack_1, ack => sendB_CP_2093_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	52 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/ptr_deref_956_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/ptr_deref_956_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/ptr_deref_956_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/ptr_deref_956_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/word_access_start/word_0/rr
      -- 
    rr_2703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(63), ack => ptr_deref_956_store_0_req_0); -- 
    sendB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(52) & sendB_CP_2093_elements(62);
      gj_sendB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	91 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Sample/word_access_start/word_0/ra
      -- 
    ra_2704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_956_store_0_ack_0, ack => sendB_CP_2093_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	52 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	96 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_Update/word_access_complete/word_0/ca
      -- 
    ca_2715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_956_store_0_ack_1, ack => sendB_CP_2093_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_Sample/ra
      -- 
    ra_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_0, ack => sendB_CP_2093_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	52 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_967_Update/ca
      -- 
    ca_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_967_inst_ack_1, ack => sendB_CP_2093_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: 	91 
    -- CP-element group 68: 	52 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (9) 
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/ptr_deref_977_Split/$entry
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/ptr_deref_977_Split/$exit
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/ptr_deref_977_Split/split_req
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/ptr_deref_977_Split/split_ack
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/word_access_start/$entry
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/word_access_start/word_0/$entry
      -- CP-element group 68: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/word_access_start/word_0/rr
      -- 
    rr_2767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(68), ack => ptr_deref_977_store_0_req_0); -- 
    sendB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(67) & sendB_CP_2093_elements(91) & sendB_CP_2093_elements(52);
      gj_sendB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	92 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/word_access_start/$exit
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/word_access_start/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Sample/word_access_start/word_0/ra
      -- 
    ra_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_977_store_0_ack_0, ack => sendB_CP_2093_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	52 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	96 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Update/word_access_complete/$exit
      -- CP-element group 70: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Update/word_access_complete/word_0/$exit
      -- CP-element group 70: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_Update/word_access_complete/word_0/ca
      -- 
    ca_2779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_977_store_0_ack_1, ack => sendB_CP_2093_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	60 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_Sample/ra
      -- 
    ra_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_988_inst_ack_0, ack => sendB_CP_2093_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	52 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_988_Update/ca
      -- 
    ca_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_988_inst_ack_1, ack => sendB_CP_2093_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: 	92 
    -- CP-element group 73: 	52 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (9) 
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/ptr_deref_998_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/ptr_deref_998_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/ptr_deref_998_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/ptr_deref_998_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_sample_start_
      -- 
    rr_2831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(73), ack => ptr_deref_998_store_0_req_0); -- 
    sendB_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(72) & sendB_CP_2093_elements(92) & sendB_CP_2093_elements(52);
      gj_sendB_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	93 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/word_access_start/word_0/ra
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_sample_completed_
      -- 
    ra_2832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_998_store_0_ack_0, ack => sendB_CP_2093_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	52 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	96 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_Update/word_access_complete/word_0/ca
      -- 
    ca_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_998_store_0_ack_1, ack => sendB_CP_2093_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	60 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_sample_completed_
      -- 
    ra_2852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1009_inst_ack_0, ack => sendB_CP_2093_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	52 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1009_update_completed_
      -- 
    ca_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1009_inst_ack_1, ack => sendB_CP_2093_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: 	93 
    -- CP-element group 78: 	52 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/ptr_deref_1019_Split/split_ack
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/word_access_start/$entry
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/word_access_start/word_0/$entry
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/word_access_start/word_0/rr
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/ptr_deref_1019_Split/split_req
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/ptr_deref_1019_Split/$exit
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/ptr_deref_1019_Split/$entry
      -- CP-element group 78: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/$entry
      -- 
    rr_2895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(78), ack => ptr_deref_1019_store_0_req_0); -- 
    sendB_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(77) & sendB_CP_2093_elements(93) & sendB_CP_2093_elements(52);
      gj_sendB_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	94 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/word_access_start/$exit
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/word_access_start/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/word_access_start/word_0/ra
      -- CP-element group 79: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Sample/$exit
      -- 
    ra_2896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1019_store_0_ack_0, ack => sendB_CP_2093_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	52 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	96 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Update/word_access_complete/$exit
      -- CP-element group 80: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Update/word_access_complete/word_0/ca
      -- CP-element group 80: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Update/word_access_complete/word_0/$exit
      -- CP-element group 80: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_Update/$exit
      -- 
    ca_2907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1019_store_0_ack_1, ack => sendB_CP_2093_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	60 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_sample_completed_
      -- 
    ra_2916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1030_inst_ack_0, ack => sendB_CP_2093_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	52 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1030_update_completed_
      -- 
    ca_2921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1030_inst_ack_1, ack => sendB_CP_2093_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: 	94 
    -- CP-element group 83: 	52 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/ptr_deref_1040_Split/$entry
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/ptr_deref_1040_Split/$exit
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/ptr_deref_1040_Split/split_req
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/ptr_deref_1040_Split/split_ack
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/word_access_start/$entry
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/word_access_start/word_0/$entry
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/word_access_start/word_0/rr
      -- CP-element group 83: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_sample_start_
      -- 
    rr_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(83), ack => ptr_deref_1040_store_0_req_0); -- 
    sendB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(82) & sendB_CP_2093_elements(94) & sendB_CP_2093_elements(52);
      gj_sendB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	95 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/word_access_start/$exit
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/word_access_start/word_0/$exit
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Sample/word_access_start/word_0/ra
      -- CP-element group 84: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_sample_completed_
      -- 
    ra_2960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1040_store_0_ack_0, ack => sendB_CP_2093_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	52 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	96 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Update/word_access_complete/word_0/ca
      -- CP-element group 85: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Update/word_access_complete/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Update/word_access_complete/$exit
      -- CP-element group 85: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_Update/$exit
      -- 
    ca_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1040_store_0_ack_1, ack => sendB_CP_2093_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	60 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_sample_completed_
      -- 
    ra_2980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1051_inst_ack_0, ack => sendB_CP_2093_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	52 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/type_cast_1051_update_completed_
      -- 
    ca_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1051_inst_ack_1, ack => sendB_CP_2093_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: 	95 
    -- CP-element group 88: 	52 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/ptr_deref_1061_Split/split_req
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/ptr_deref_1061_Split/split_ack
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/word_access_start/$entry
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/word_access_start/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/word_access_start/word_0/rr
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/ptr_deref_1061_Split/$exit
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/ptr_deref_1061_Split/$entry
      -- CP-element group 88: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/$entry
      -- 
    rr_3023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(88), ack => ptr_deref_1061_store_0_req_0); -- 
    sendB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(87) & sendB_CP_2093_elements(95) & sendB_CP_2093_elements(52);
      gj_sendB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/word_access_start/$exit
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/word_access_start/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/word_access_start/word_0/ra
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Sample/$exit
      -- 
    ra_3024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1061_store_0_ack_0, ack => sendB_CP_2093_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	52 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	96 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Update/word_access_complete/word_0/ca
      -- CP-element group 90: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Update/word_access_complete/word_0/$exit
      -- CP-element group 90: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1061_Update/word_access_complete/$exit
      -- 
    ca_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1061_store_0_ack_1, ack => sendB_CP_2093_elements(90)); -- 
    -- CP-element group 91:  transition  delay-element  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	64 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	68 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_956_ptr_deref_977_delay
      -- 
    -- Element group sendB_CP_2093_elements(91) is a control-delay.
    cp_element_91_delay: control_delay_element  generic map(name => " 91_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(64), ack => sendB_CP_2093_elements(91), clk => clk, reset =>reset);
    -- CP-element group 92:  transition  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	69 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	73 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_977_ptr_deref_998_delay
      -- 
    -- Element group sendB_CP_2093_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(69), ack => sendB_CP_2093_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  transition  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	74 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	78 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_998_ptr_deref_1019_delay
      -- 
    -- Element group sendB_CP_2093_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(74), ack => sendB_CP_2093_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  transition  delay-element  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	79 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	83 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1019_ptr_deref_1040_delay
      -- 
    -- Element group sendB_CP_2093_elements(94) is a control-delay.
    cp_element_94_delay: control_delay_element  generic map(name => " 94_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(79), ack => sendB_CP_2093_elements(94), clk => clk, reset =>reset);
    -- CP-element group 95:  transition  delay-element  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	84 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	88 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/ptr_deref_1040_ptr_deref_1061_delay
      -- 
    -- Element group sendB_CP_2093_elements(95) is a control-delay.
    cp_element_95_delay: control_delay_element  generic map(name => " 95_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(84), ack => sendB_CP_2093_elements(95), clk => clk, reset =>reset);
    -- CP-element group 96:  branch  join  transition  place  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	70 
    -- CP-element group 96: 	65 
    -- CP-element group 96: 	75 
    -- CP-element group 96: 	80 
    -- CP-element group 96: 	85 
    -- CP-element group 96: 	90 
    -- CP-element group 96: 	54 
    -- CP-element group 96: 	55 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (10) 
      -- CP-element group 96: 	 branch_block_stmt_689/if_stmt_1070__entry__
      -- CP-element group 96: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069__exit__
      -- CP-element group 96: 	 branch_block_stmt_689/assign_stmt_926_to_assign_stmt_1069/$exit
      -- CP-element group 96: 	 branch_block_stmt_689/if_stmt_1070_else_link/$entry
      -- CP-element group 96: 	 branch_block_stmt_689/if_stmt_1070_if_link/$entry
      -- CP-element group 96: 	 branch_block_stmt_689/if_stmt_1070_eval_test/branch_req
      -- CP-element group 96: 	 branch_block_stmt_689/if_stmt_1070_eval_test/$exit
      -- CP-element group 96: 	 branch_block_stmt_689/if_stmt_1070_eval_test/$entry
      -- CP-element group 96: 	 branch_block_stmt_689/R_cmp53x_xi_1071_place
      -- CP-element group 96: 	 branch_block_stmt_689/if_stmt_1070_dead_link/$entry
      -- 
    branch_req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(96), ack => if_stmt_1070_branch_req_0); -- 
    sendB_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(70) & sendB_CP_2093_elements(65) & sendB_CP_2093_elements(75) & sendB_CP_2093_elements(80) & sendB_CP_2093_elements(85) & sendB_CP_2093_elements(90) & sendB_CP_2093_elements(54) & sendB_CP_2093_elements(55);
      gj_sendB_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  place  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	137 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_689/ifx_xthen_sendRemainingElementsx_xexit
      -- CP-element group 97: 	 branch_block_stmt_689/if_stmt_1070_if_link/if_choice_transition
      -- CP-element group 97: 	 branch_block_stmt_689/if_stmt_1070_if_link/$exit
      -- CP-element group 97: 	 branch_block_stmt_689/ifx_xthen_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 97: 	 branch_block_stmt_689/ifx_xthen_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1070_branch_ack_1, ack => sendB_CP_2093_elements(97)); -- 
    -- CP-element group 98:  merge  transition  place  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	131 
    -- CP-element group 98:  members (18) 
      -- CP-element group 98: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_1082_to_assign_stmt_1107__entry__
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_1082_to_assign_stmt_1107__exit__
      -- CP-element group 98: 	 branch_block_stmt_689/merge_stmt_1076__exit__
      -- CP-element group 98: 	 branch_block_stmt_689/ifx_xthen_bbx_xnphx_xi
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_1082_to_assign_stmt_1107/$exit
      -- CP-element group 98: 	 branch_block_stmt_689/assign_stmt_1082_to_assign_stmt_1107/$entry
      -- CP-element group 98: 	 branch_block_stmt_689/if_stmt_1070_else_link/else_choice_transition
      -- CP-element group 98: 	 branch_block_stmt_689/if_stmt_1070_else_link/$exit
      -- CP-element group 98: 	 branch_block_stmt_689/ifx_xthen_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 98: 	 branch_block_stmt_689/ifx_xthen_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 98: 	 branch_block_stmt_689/merge_stmt_1076_PhiReqMerge
      -- CP-element group 98: 	 branch_block_stmt_689/merge_stmt_1076_PhiAck/$entry
      -- CP-element group 98: 	 branch_block_stmt_689/merge_stmt_1076_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_689/merge_stmt_1076_PhiAck/dummy
      -- CP-element group 98: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 98: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/$entry
      -- CP-element group 98: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/$entry
      -- 
    else_choice_transition_3057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1070_branch_ack_0, ack => sendB_CP_2093_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	136 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	116 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_sample_complete
      -- 
    ack_3092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1128_index_offset_ack_0, ack => sendB_CP_2093_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	136 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (11) 
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_request/$entry
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_request/req
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_root_address_calculated
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_offset_calculated
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_base_plus_offset/sum_rename_ack
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_base_plus_offset/sum_rename_req
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_base_plus_offset/$exit
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_base_plus_offset/$entry
      -- CP-element group 100: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_Update/ack
      -- 
    ack_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1128_index_offset_ack_1, ack => sendB_CP_2093_elements(100)); -- 
    req_3106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(100), ack => array_obj_ref_1128_final_reg_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_request/$exit
      -- CP-element group 101: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_request/ack
      -- 
    ack_3107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1128_final_reg_ack_0, ack => sendB_CP_2093_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	136 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	107 
    -- CP-element group 102:  members (24) 
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_plus_offset/$entry
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_plus_offset/$exit
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_plus_offset/sum_rename_req
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_plus_offset/sum_rename_ack
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_word_addrgen/$entry
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_word_addrgen/$exit
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_word_addrgen/root_register_req
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_word_addrgen/root_register_ack
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Sample/word_access_start/$entry
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Sample/word_access_start/word_0/rr
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Sample/word_access_start/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_addr_resize/base_resize_ack
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_addr_resize/base_resize_req
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_addr_resize/$exit
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_addr_resize/$entry
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_address_resized
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_root_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_complete/ack
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_word_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_base_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_complete/$exit
      -- 
    ack_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1128_final_reg_ack_1, ack => sendB_CP_2093_elements(102)); -- 
    rr_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(102), ack => ptr_deref_1144_load_0_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	136 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	116 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_sample_complete
      -- CP-element group 103: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_Sample/ack
      -- 
    ack_3139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1140_index_offset_ack_0, ack => sendB_CP_2093_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	136 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (11) 
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_request/req
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_request/$entry
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_offset_calculated
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_base_plus_offset/sum_rename_ack
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_base_plus_offset/sum_rename_req
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_root_address_calculated
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_base_plus_offset/$exit
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_base_plus_offset/$entry
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_Update/$exit
      -- 
    ack_3144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1140_index_offset_ack_1, ack => sendB_CP_2093_elements(104)); -- 
    req_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(104), ack => array_obj_ref_1140_final_reg_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_request/ack
      -- CP-element group 105: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_request/$exit
      -- CP-element group 105: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_sample_completed_
      -- 
    ack_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1140_final_reg_ack_0, ack => sendB_CP_2093_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	136 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	111 
    -- CP-element group 106:  members (24) 
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_complete/$exit
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_complete/ack
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_addr_resize/$exit
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Sample/word_access_start/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_word_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_root_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_address_resized
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_addr_resize/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_addr_resize/base_resize_req
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_addr_resize/base_resize_ack
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_word_addrgen/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_word_addrgen/$exit
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_plus_offset/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_plus_offset/$exit
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Sample/word_access_start/word_0/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_word_addrgen/root_register_req
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_plus_offset/sum_rename_req
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_plus_offset/sum_rename_ack
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_word_addrgen/root_register_ack
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_base_address_calculated
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Sample/word_access_start/word_0/rr
      -- 
    ack_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1140_final_reg_ack_1, ack => sendB_CP_2093_elements(106)); -- 
    rr_3256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(106), ack => ptr_deref_1151_load_0_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	102 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Sample/word_access_start/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Sample/word_access_start/$exit
      -- CP-element group 107: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Sample/word_access_start/word_0/ra
      -- 
    ra_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1144_load_0_ack_0, ack => sendB_CP_2093_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	136 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (12) 
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_Sample/req
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/word_access_complete/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/ptr_deref_1144_Merge/merge_req
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/ptr_deref_1144_Merge/$entry
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/ptr_deref_1144_Merge/$exit
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/word_access_complete/$exit
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/word_access_complete/word_0/ca
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/ptr_deref_1144_Merge/merge_ack
      -- CP-element group 108: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_Sample/$entry
      -- 
    ca_3204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1144_load_0_ack_1, ack => sendB_CP_2093_elements(108)); -- 
    req_3217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(108), ack => WPIPE_maxpool_output_pipe_1146_inst_req_0); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_update_start_
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_Sample/ack
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_Update/req
      -- CP-element group 109: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_Sample/$exit
      -- 
    ack_3218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1146_inst_ack_0, ack => sendB_CP_2093_elements(109)); -- 
    req_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(109), ack => WPIPE_maxpool_output_pipe_1146_inst_req_1); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	113 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_Update/ack
      -- CP-element group 110: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1146_Update/$exit
      -- 
    ack_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1146_inst_ack_1, ack => sendB_CP_2093_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	106 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Sample/word_access_start/$exit
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Sample/word_access_start/word_0/ra
      -- CP-element group 111: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Sample/word_access_start/word_0/$exit
      -- 
    ra_3257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1151_load_0_ack_0, ack => sendB_CP_2093_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	136 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/word_access_complete/$exit
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/word_access_complete/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/ptr_deref_1151_Merge/$exit
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/ptr_deref_1151_Merge/merge_req
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/word_access_complete/word_0/ca
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/ptr_deref_1151_Merge/$entry
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/ptr_deref_1151_Merge/merge_ack
      -- 
    ca_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1151_load_0_ack_1, ack => sendB_CP_2093_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	110 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_Sample/req
      -- 
    req_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(113), ack => WPIPE_maxpool_output_pipe_1153_inst_req_0); -- 
    sendB_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(110) & sendB_CP_2093_elements(112);
      gj_sendB_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_update_start_
      -- CP-element group 114: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_Update/req
      -- 
    ack_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1153_inst_ack_0, ack => sendB_CP_2093_elements(114)); -- 
    req_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(114), ack => WPIPE_maxpool_output_pipe_1153_inst_req_1); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/WPIPE_maxpool_output_pipe_1153_Update/ack
      -- 
    ack_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1153_inst_ack_1, ack => sendB_CP_2093_elements(115)); -- 
    -- CP-element group 116:  branch  join  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	99 
    -- CP-element group 116: 	103 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_689/if_stmt_1167__entry__
      -- CP-element group 116: 	 branch_block_stmt_689/R_exitcond1_1168_place
      -- CP-element group 116: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166__exit__
      -- CP-element group 116: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/$exit
      -- CP-element group 116: 	 branch_block_stmt_689/if_stmt_1167_dead_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_689/if_stmt_1167_eval_test/$entry
      -- CP-element group 116: 	 branch_block_stmt_689/if_stmt_1167_eval_test/$exit
      -- CP-element group 116: 	 branch_block_stmt_689/if_stmt_1167_eval_test/branch_req
      -- CP-element group 116: 	 branch_block_stmt_689/if_stmt_1167_if_link/$entry
      -- CP-element group 116: 	 branch_block_stmt_689/if_stmt_1167_else_link/$entry
      -- 
    branch_req_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(116), ack => if_stmt_1167_branch_req_0); -- 
    sendB_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(99) & sendB_CP_2093_elements(103) & sendB_CP_2093_elements(115);
      gj_sendB_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  merge  transition  place  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	137 
    -- CP-element group 117:  members (13) 
      -- CP-element group 117: 	 branch_block_stmt_689/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit
      -- CP-element group 117: 	 branch_block_stmt_689/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit
      -- CP-element group 117: 	 branch_block_stmt_689/merge_stmt_1173__exit__
      -- CP-element group 117: 	 branch_block_stmt_689/if_stmt_1167_if_link/$exit
      -- CP-element group 117: 	 branch_block_stmt_689/if_stmt_1167_if_link/if_choice_transition
      -- CP-element group 117: 	 branch_block_stmt_689/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit_PhiReq/$entry
      -- CP-element group 117: 	 branch_block_stmt_689/forx_xbodyx_xi_sendRemainingElementsx_xexitx_xloopexit_PhiReq/$exit
      -- CP-element group 117: 	 branch_block_stmt_689/merge_stmt_1173_PhiReqMerge
      -- CP-element group 117: 	 branch_block_stmt_689/merge_stmt_1173_PhiAck/$entry
      -- CP-element group 117: 	 branch_block_stmt_689/merge_stmt_1173_PhiAck/$exit
      -- CP-element group 117: 	 branch_block_stmt_689/merge_stmt_1173_PhiAck/dummy
      -- CP-element group 117: 	 branch_block_stmt_689/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 117: 	 branch_block_stmt_689/sendRemainingElementsx_xexitx_xloopexit_sendRemainingElementsx_xexit_PhiReq/$exit
      -- 
    if_choice_transition_3300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1167_branch_ack_1, ack => sendB_CP_2093_elements(117)); -- 
    -- CP-element group 118:  fork  transition  place  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	132 
    -- CP-element group 118: 	133 
    -- CP-element group 118:  members (12) 
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 118: 	 branch_block_stmt_689/if_stmt_1167_else_link/$exit
      -- CP-element group 118: 	 branch_block_stmt_689/if_stmt_1167_else_link/else_choice_transition
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/$entry
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/$entry
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/$entry
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/$entry
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1167_branch_ack_0, ack => sendB_CP_2093_elements(118)); -- 
    rr_3468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(118), ack => type_cast_1116_inst_req_0); -- 
    cr_3473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(118), ack => type_cast_1116_inst_req_1); -- 
    -- CP-element group 119:  transition  output  delay-element  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	1 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_689/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_689/bbx_xnph_forx_xbody_PhiReq/phi_stmt_736/$exit
      -- CP-element group 119: 	 branch_block_stmt_689/bbx_xnph_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_689/bbx_xnph_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_740_konst_delay_trans
      -- CP-element group 119: 	 branch_block_stmt_689/bbx_xnph_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_req
      -- 
    phi_stmt_736_req_3329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_736_req_3329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(119), ack => phi_stmt_736_req_0); -- 
    -- Element group sendB_CP_2093_elements(119) is a control-delay.
    cp_element_119_delay: control_delay_element  generic map(name => " 119_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(1), ack => sendB_CP_2093_elements(119), clk => clk, reset =>reset);
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	50 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/Sample/ra
      -- 
    ra_3349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_742_inst_ack_0, ack => sendB_CP_2093_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	50 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/Update/ca
      -- 
    ca_3354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_742_inst_ack_1, ack => sendB_CP_2093_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (6) 
      -- CP-element group 122: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/$exit
      -- CP-element group 122: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/$exit
      -- CP-element group 122: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/$exit
      -- CP-element group 122: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_sources/type_cast_742/SplitProtocol/$exit
      -- CP-element group 122: 	 branch_block_stmt_689/forx_xbody_forx_xbody_PhiReq/phi_stmt_736/phi_stmt_736_req
      -- 
    phi_stmt_736_req_3355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_736_req_3355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(122), ack => phi_stmt_736_req_1); -- 
    sendB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(120) & sendB_CP_2093_elements(121);
      gj_sendB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_689/merge_stmt_735_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_689/merge_stmt_735_PhiAck/$entry
      -- 
    sendB_CP_2093_elements(123) <= OrReduce(sendB_CP_2093_elements(119) & sendB_CP_2093_elements(122));
    -- CP-element group 124:  fork  transition  place  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	6 
    -- CP-element group 124: 	8 
    -- CP-element group 124: 	10 
    -- CP-element group 124: 	12 
    -- CP-element group 124: 	14 
    -- CP-element group 124: 	16 
    -- CP-element group 124: 	18 
    -- CP-element group 124: 	20 
    -- CP-element group 124: 	22 
    -- CP-element group 124: 	24 
    -- CP-element group 124: 	3 
    -- CP-element group 124: 	4 
    -- CP-element group 124:  members (53) 
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_scaled_1
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_resized_1
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_Update/req
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_Sample/req
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_scale_1/scale_rename_req
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_resize_1/$exit
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_resize_1/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_resize_1/index_resize_req
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_scale_1/scale_rename_ack
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863__entry__
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_update_start
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_resize_1/index_resize_ack
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_scale_1/$exit
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_scale_1/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_final_index_sum_regn_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/array_obj_ref_748_index_computed_1
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/merge_stmt_735__exit__
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_complete/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/addr_of_749_complete/req
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/word_access_complete/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/word_access_complete/word_0/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/ptr_deref_753_Update/word_access_complete/word_0/cr
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_757_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_767_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_777_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_787_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_797_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_807_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_817_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_update_start_
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_689/assign_stmt_750_to_assign_stmt_863/type_cast_827_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_689/merge_stmt_735_PhiAck/$exit
      -- CP-element group 124: 	 branch_block_stmt_689/merge_stmt_735_PhiAck/phi_stmt_736_ack
      -- 
    phi_stmt_736_ack_3360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_736_ack_0, ack => sendB_CP_2093_elements(124)); -- 
    req_2204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => array_obj_ref_748_index_offset_req_1); -- 
    req_2199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => array_obj_ref_748_index_offset_req_0); -- 
    req_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => addr_of_749_final_reg_req_1); -- 
    cr_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => ptr_deref_753_load_0_req_1); -- 
    cr_2283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => type_cast_757_inst_req_1); -- 
    cr_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => type_cast_767_inst_req_1); -- 
    cr_2311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => type_cast_777_inst_req_1); -- 
    cr_2325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => type_cast_787_inst_req_1); -- 
    cr_2339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => type_cast_797_inst_req_1); -- 
    cr_2353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => type_cast_807_inst_req_1); -- 
    cr_2367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => type_cast_817_inst_req_1); -- 
    cr_2381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(124), ack => type_cast_827_inst_req_1); -- 
    -- CP-element group 125:  transition  output  delay-element  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	2 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	129 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/$exit
      -- CP-element group 125: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_896/$exit
      -- CP-element group 125: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/$exit
      -- CP-element group 125: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_902_konst_delay_trans
      -- CP-element group 125: 	 branch_block_stmt_689/entry_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_req
      -- 
    phi_stmt_896_req_3383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_896_req_3383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(125), ack => phi_stmt_896_req_1); -- 
    -- Element group sendB_CP_2093_elements(125) is a control-delay.
    cp_element_125_delay: control_delay_element  generic map(name => " 125_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(2), ack => sendB_CP_2093_elements(125), clk => clk, reset =>reset);
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	49 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/Sample/ra
      -- 
    ra_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_899_inst_ack_0, ack => sendB_CP_2093_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	49 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/Update/ca
      -- 
    ca_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_899_inst_ack_1, ack => sendB_CP_2093_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 128: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/$exit
      -- CP-element group 128: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/$exit
      -- CP-element group 128: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/$exit
      -- CP-element group 128: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_sources/type_cast_899/SplitProtocol/$exit
      -- CP-element group 128: 	 branch_block_stmt_689/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_896/phi_stmt_896_req
      -- 
    phi_stmt_896_req_3409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_896_req_3409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(128), ack => phi_stmt_896_req_0); -- 
    sendB_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(126) & sendB_CP_2093_elements(127);
      gj_sendB_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  merge  transition  place  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	125 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_689/merge_stmt_895_PhiReqMerge
      -- CP-element group 129: 	 branch_block_stmt_689/merge_stmt_895_PhiAck/$entry
      -- 
    sendB_CP_2093_elements(129) <= OrReduce(sendB_CP_2093_elements(125) & sendB_CP_2093_elements(128));
    -- CP-element group 130:  branch  transition  place  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	51 
    -- CP-element group 130: 	52 
    -- CP-element group 130:  members (15) 
      -- CP-element group 130: 	 branch_block_stmt_689/assign_stmt_909_to_assign_stmt_915__entry__
      -- CP-element group 130: 	 branch_block_stmt_689/if_stmt_916__entry__
      -- CP-element group 130: 	 branch_block_stmt_689/assign_stmt_909_to_assign_stmt_915__exit__
      -- CP-element group 130: 	 branch_block_stmt_689/merge_stmt_895__exit__
      -- CP-element group 130: 	 branch_block_stmt_689/assign_stmt_909_to_assign_stmt_915/$entry
      -- CP-element group 130: 	 branch_block_stmt_689/assign_stmt_909_to_assign_stmt_915/$exit
      -- CP-element group 130: 	 branch_block_stmt_689/if_stmt_916_dead_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_689/if_stmt_916_eval_test/$entry
      -- CP-element group 130: 	 branch_block_stmt_689/if_stmt_916_eval_test/$exit
      -- CP-element group 130: 	 branch_block_stmt_689/if_stmt_916_eval_test/branch_req
      -- CP-element group 130: 	 branch_block_stmt_689/R_tobool_917_place
      -- CP-element group 130: 	 branch_block_stmt_689/if_stmt_916_if_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_689/if_stmt_916_else_link/$entry
      -- CP-element group 130: 	 branch_block_stmt_689/merge_stmt_895_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_689/merge_stmt_895_PhiAck/phi_stmt_896_ack
      -- 
    phi_stmt_896_ack_3414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_896_ack_0, ack => sendB_CP_2093_elements(130)); -- 
    branch_req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(130), ack => if_stmt_916_branch_req_0); -- 
    -- CP-element group 131:  transition  output  delay-element  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	98 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	135 
    -- CP-element group 131:  members (5) 
      -- CP-element group 131: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- CP-element group 131: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/$exit
      -- CP-element group 131: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/$exit
      -- CP-element group 131: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1114_konst_delay_trans
      -- CP-element group 131: 	 branch_block_stmt_689/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_req
      -- 
    phi_stmt_1110_req_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1110_req_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(131), ack => phi_stmt_1110_req_0); -- 
    -- Element group sendB_CP_2093_elements(131) is a control-delay.
    cp_element_131_delay: control_delay_element  generic map(name => " 131_delay", delay_value => 1)  port map(req => sendB_CP_2093_elements(98), ack => sendB_CP_2093_elements(131), clk => clk, reset =>reset);
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	118 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/Sample/ra
      -- 
    ra_3469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1116_inst_ack_0, ack => sendB_CP_2093_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	118 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (2) 
      -- CP-element group 133: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/Update/ca
      -- 
    ca_3474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1116_inst_ack_1, ack => sendB_CP_2093_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- CP-element group 134: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/$exit
      -- CP-element group 134: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/$exit
      -- CP-element group 134: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/$exit
      -- CP-element group 134: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_sources/type_cast_1116/SplitProtocol/$exit
      -- CP-element group 134: 	 branch_block_stmt_689/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1110/phi_stmt_1110_req
      -- 
    phi_stmt_1110_req_3475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1110_req_3475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(134), ack => phi_stmt_1110_req_1); -- 
    sendB_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "sendB_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2093_elements(132) & sendB_CP_2093_elements(133);
      gj_sendB_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2093_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  merge  transition  place  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	131 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_689/merge_stmt_1109_PhiReqMerge
      -- CP-element group 135: 	 branch_block_stmt_689/merge_stmt_1109_PhiAck/$entry
      -- 
    sendB_CP_2093_elements(135) <= OrReduce(sendB_CP_2093_elements(131) & sendB_CP_2093_elements(134));
    -- CP-element group 136:  fork  transition  place  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	99 
    -- CP-element group 136: 	100 
    -- CP-element group 136: 	102 
    -- CP-element group 136: 	103 
    -- CP-element group 136: 	104 
    -- CP-element group 136: 	106 
    -- CP-element group 136: 	108 
    -- CP-element group 136: 	112 
    -- CP-element group 136:  members (53) 
      -- CP-element group 136: 	 branch_block_stmt_689/merge_stmt_1109__exit__
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166__entry__
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_scale_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_update_start_
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_scale_1/scale_rename_req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_computed_1
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_resize_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_scale_1/scale_rename_ack
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_resize_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_resize_1/index_resize_req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_resize_1/index_resize_ack
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_resized_1
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_scale_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_scale_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_scale_1/scale_rename_req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_complete/req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/word_access_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_scale_1/scale_rename_ack
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_Sample/req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_update_start
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_scaled_1
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/word_access_complete/word_0/cr
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_Update/word_access_complete/word_0/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/word_access_complete/word_0/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1151_update_start_
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_update_start
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_update_start_
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/word_access_complete/word_0/cr
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_final_index_sum_regn_Update/req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_Sample/req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/word_access_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_computed_1
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_scaled_1
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_scale_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_resize_1/index_resize_ack
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_index_resized_1
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/ptr_deref_1144_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_update_start_
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_resize_1/index_resize_req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_resize_1/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_index_resize_1/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_complete/req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1140_final_index_sum_regn_Update/req
      -- CP-element group 136: 	 branch_block_stmt_689/assign_stmt_1123_to_assign_stmt_1166/array_obj_ref_1128_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_689/merge_stmt_1109_PhiAck/$exit
      -- CP-element group 136: 	 branch_block_stmt_689/merge_stmt_1109_PhiAck/phi_stmt_1110_ack
      -- 
    phi_stmt_1110_ack_3480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1110_ack_0, ack => sendB_CP_2093_elements(136)); -- 
    req_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => array_obj_ref_1140_final_reg_req_1); -- 
    req_3091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => array_obj_ref_1128_index_offset_req_0); -- 
    cr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => ptr_deref_1151_load_0_req_1); -- 
    cr_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => ptr_deref_1144_load_0_req_1); -- 
    req_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => array_obj_ref_1128_index_offset_req_1); -- 
    req_3138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => array_obj_ref_1140_index_offset_req_0); -- 
    req_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => array_obj_ref_1128_final_reg_req_1); -- 
    req_3143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2093_elements(136), ack => array_obj_ref_1140_index_offset_req_1); -- 
    -- CP-element group 137:  merge  transition  place  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	97 
    -- CP-element group 137: 	117 
    -- CP-element group 137: 	51 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (16) 
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1177__exit__
      -- CP-element group 137: 	 branch_block_stmt_689/return__
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1175__exit__
      -- CP-element group 137: 	 $exit
      -- CP-element group 137: 	 branch_block_stmt_689/$exit
      -- CP-element group 137: 	 branch_block_stmt_689/branch_block_stmt_689__exit__
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1177_PhiReqMerge
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1175_PhiReqMerge
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1175_PhiAck/$entry
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1175_PhiAck/$exit
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1175_PhiAck/dummy
      -- CP-element group 137: 	 branch_block_stmt_689/return___PhiReq/$entry
      -- CP-element group 137: 	 branch_block_stmt_689/return___PhiReq/$exit
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1177_PhiAck/$entry
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1177_PhiAck/$exit
      -- CP-element group 137: 	 branch_block_stmt_689/merge_stmt_1177_PhiAck/dummy
      -- 
    sendB_CP_2093_elements(137) <= OrReduce(sendB_CP_2093_elements(97) & sendB_CP_2093_elements(117) & sendB_CP_2093_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_891_wire : std_logic_vector(63 downto 0);
    signal R_indvar_747_resized : std_logic_vector(13 downto 0);
    signal R_indvar_747_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_930_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_930_scaled : std_logic_vector(13 downto 0);
    signal R_tmp2_1127_resized : std_logic_vector(2 downto 0);
    signal R_tmp2_1127_scaled : std_logic_vector(2 downto 0);
    signal R_tmp3_1139_resized : std_logic_vector(2 downto 0);
    signal R_tmp3_1139_scaled : std_logic_vector(2 downto 0);
    signal and70_909 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1128_constant_part_of_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1128_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1128_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1128_offset_scale_factor_1 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1128_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1128_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1140_constant_part_of_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1140_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1140_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1140_offset_scale_factor_1 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1140_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1140_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_748_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_748_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_748_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_748_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_748_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_748_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_931_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_931_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_931_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_931_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_931_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_931_root_address : std_logic_vector(13 downto 0);
    signal arrayidx11x_xi_975 : std_logic_vector(31 downto 0);
    signal arrayidx17x_xi_996 : std_logic_vector(31 downto 0);
    signal arrayidx23x_xi_1017 : std_logic_vector(31 downto 0);
    signal arrayidx29x_xi_1038 : std_logic_vector(31 downto 0);
    signal arrayidx35x_xi_1059 : std_logic_vector(31 downto 0);
    signal arrayidx43x_xi_1129 : std_logic_vector(31 downto 0);
    signal arrayidx48x_xi_1141 : std_logic_vector(31 downto 0);
    signal arrayidx5x_xi_954 : std_logic_vector(31 downto 0);
    signal arrayidx_750 : std_logic_vector(31 downto 0);
    signal arrayidxx_xi_933 : std_logic_vector(31 downto 0);
    signal cmp53x_xi_1069 : std_logic_vector(0 downto 0);
    signal cmp77_701 : std_logic_vector(0 downto 0);
    signal conv10x_xi_968 : std_logic_vector(7 downto 0);
    signal conv14_768 : std_logic_vector(7 downto 0);
    signal conv16x_xi_989 : std_logic_vector(7 downto 0);
    signal conv20_778 : std_logic_vector(7 downto 0);
    signal conv22x_xi_1010 : std_logic_vector(7 downto 0);
    signal conv26_788 : std_logic_vector(7 downto 0);
    signal conv28x_xi_1031 : std_logic_vector(7 downto 0);
    signal conv32_798 : std_logic_vector(7 downto 0);
    signal conv34x_xi_1052 : std_logic_vector(7 downto 0);
    signal conv38_808 : std_logic_vector(7 downto 0);
    signal conv44_818 : std_logic_vector(7 downto 0);
    signal conv50_828 : std_logic_vector(7 downto 0);
    signal conv74_926 : std_logic_vector(15 downto 0);
    signal conv8_758 : std_logic_vector(7 downto 0);
    signal convx_xi_947 : std_logic_vector(7 downto 0);
    signal exitcond1_1166 : std_logic_vector(0 downto 0);
    signal exitcond_863 : std_logic_vector(0 downto 0);
    signal iNsTr_29_1094 : std_logic_vector(63 downto 0);
    signal indvar_736 : std_logic_vector(63 downto 0);
    signal indvarx_xi_1110 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_858 : std_logic_vector(63 downto 0);
    signal indvarx_xnextx_xi_1161 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_896 : std_logic_vector(63 downto 0);
    signal out_datax_xi_695 : std_logic_vector(31 downto 0);
    signal phitmp_893 : std_logic_vector(63 downto 0);
    signal ptr_deref_1019_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1019_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1019_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1019_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1019_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1019_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1040_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1040_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1040_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1040_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1040_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1040_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1061_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1061_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1061_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1061_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1061_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1061_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1144_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1144_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1144_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1144_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1144_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1151_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1151_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1151_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1151_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1151_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_753_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_753_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_753_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_753_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_753_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_936_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_936_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_936_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_936_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_936_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_956_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_956_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_956_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_956_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_956_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_956_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_977_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_977_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_977_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_977_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_977_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_977_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_998_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_998_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_998_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_998_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_998_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_998_word_offset_0 : std_logic_vector(2 downto 0);
    signal shr11_764 : std_logic_vector(63 downto 0);
    signal shr13x_xi_985 : std_logic_vector(63 downto 0);
    signal shr17_774 : std_logic_vector(63 downto 0);
    signal shr19x_xi_1006 : std_logic_vector(63 downto 0);
    signal shr23_784 : std_logic_vector(63 downto 0);
    signal shr25x_xi_1027 : std_logic_vector(63 downto 0);
    signal shr29_794 : std_logic_vector(63 downto 0);
    signal shr31x_xi_1048 : std_logic_vector(63 downto 0);
    signal shr35_804 : std_logic_vector(63 downto 0);
    signal shr41_814 : std_logic_vector(63 downto 0);
    signal shr47_824 : std_logic_vector(63 downto 0);
    signal shr7x_xi_964 : std_logic_vector(63 downto 0);
    signal shr_714 : std_logic_vector(63 downto 0);
    signal shrx_xi_943 : std_logic_vector(63 downto 0);
    signal tmp1x_xi_937 : std_logic_vector(63 downto 0);
    signal tmp2_1123 : std_logic_vector(63 downto 0);
    signal tmp3_1135 : std_logic_vector(63 downto 0);
    signal tmp44x_xi_1145 : std_logic_vector(7 downto 0);
    signal tmp49x_xi_1152 : std_logic_vector(7 downto 0);
    signal tmp55x_xi_1082 : std_logic_vector(0 downto 0);
    signal tmp58x_xi_1107 : std_logic_vector(63 downto 0);
    signal tmp5_754 : std_logic_vector(63 downto 0);
    signal tmp80_720 : std_logic_vector(0 downto 0);
    signal tmp81_883 : std_logic_vector(63 downto 0);
    signal tmp_726 : std_logic_vector(0 downto 0);
    signal tmpx_xopx_xi_1088 : std_logic_vector(63 downto 0);
    signal tobool_915 : std_logic_vector(0 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1025_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1046_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1067_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1080_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1086_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1092_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1098_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1105_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1114_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1116_wire : std_logic_vector(63 downto 0);
    signal type_cast_1121_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1133_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1159_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_699_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_712_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_718_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_731_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_740_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_742_wire : std_logic_vector(63 downto 0);
    signal type_cast_762_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_772_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_782_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_792_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_802_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_812_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_822_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_856_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_875_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_881_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_887_wire : std_logic_vector(63 downto 0);
    signal type_cast_890_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_899_wire : std_logic_vector(63 downto 0);
    signal type_cast_902_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_907_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_913_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_941_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_962_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_983_wire_constant : std_logic_vector(63 downto 0);
    signal umax4_733 : std_logic_vector(63 downto 0);
    signal umax_877 : std_logic_vector(63 downto 0);
    signal xx_xopx_xi_1100 : std_logic_vector(63 downto 0);
    signal xxsendBxxbodyxxout_datax_xi_alloc_base_address : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    array_obj_ref_1128_constant_part_of_offset <= "000";
    array_obj_ref_1128_offset_scale_factor_0 <= "110";
    array_obj_ref_1128_offset_scale_factor_1 <= "001";
    array_obj_ref_1128_resized_base_address <= "000";
    array_obj_ref_1140_constant_part_of_offset <= "000";
    array_obj_ref_1140_offset_scale_factor_0 <= "110";
    array_obj_ref_1140_offset_scale_factor_1 <= "001";
    array_obj_ref_1140_resized_base_address <= "000";
    array_obj_ref_748_constant_part_of_offset <= "00000000000000";
    array_obj_ref_748_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_748_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_748_resized_base_address <= "00000000000000";
    array_obj_ref_931_constant_part_of_offset <= "00000000000000";
    array_obj_ref_931_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_931_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_931_resized_base_address <= "00000000000000";
    arrayidx11x_xi_975 <= "00000000000000000000000000000100";
    arrayidx17x_xi_996 <= "00000000000000000000000000000011";
    arrayidx23x_xi_1017 <= "00000000000000000000000000000010";
    arrayidx29x_xi_1038 <= "00000000000000000000000000000001";
    arrayidx35x_xi_1059 <= "00000000000000000000000000000000";
    arrayidx5x_xi_954 <= "00000000000000000000000000000101";
    out_datax_xi_695 <= "00000000000000000000000000000000";
    ptr_deref_1019_word_offset_0 <= "000";
    ptr_deref_1040_word_offset_0 <= "000";
    ptr_deref_1061_word_offset_0 <= "000";
    ptr_deref_1144_word_offset_0 <= "000";
    ptr_deref_1151_word_offset_0 <= "000";
    ptr_deref_753_word_offset_0 <= "00000000000000";
    ptr_deref_936_word_offset_0 <= "00000000000000";
    ptr_deref_956_word_offset_0 <= "000";
    ptr_deref_977_word_offset_0 <= "000";
    ptr_deref_998_word_offset_0 <= "000";
    type_cast_1004_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1025_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1046_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1067_wire_constant <= "0000000000000000";
    type_cast_1080_wire_constant <= "0000000000000001";
    type_cast_1086_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_1092_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_1098_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1105_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1114_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1121_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1133_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1159_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_699_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_712_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_718_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_724_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_731_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_740_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_762_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_772_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_782_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_792_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_802_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_812_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_822_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_856_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_875_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_881_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_890_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_902_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_907_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_913_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_941_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_962_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_983_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    xxsendBxxbodyxxout_datax_xi_alloc_base_address <= "000";
    phi_stmt_1110: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1114_wire_constant & type_cast_1116_wire;
      req <= phi_stmt_1110_req_0 & phi_stmt_1110_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1110",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1110_ack_0,
          idata => idata,
          odata => indvarx_xi_1110,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1110
    phi_stmt_736: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_740_wire_constant & type_cast_742_wire;
      req <= phi_stmt_736_req_0 & phi_stmt_736_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_736",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_736_ack_0,
          idata => idata,
          odata => indvar_736,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_736
    phi_stmt_896: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_899_wire & type_cast_902_wire_constant;
      req <= phi_stmt_896_req_0 & phi_stmt_896_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_896",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_896_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_896,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_896
    -- flow-through select operator MUX_1106_inst
    tmp58x_xi_1107 <= xx_xopx_xi_1100 when (tmp55x_xi_1082(0) /=  '0') else type_cast_1105_wire_constant;
    -- flow-through select operator MUX_732_inst
    umax4_733 <= shr_714 when (tmp_726(0) /=  '0') else type_cast_731_wire_constant;
    -- flow-through select operator MUX_876_inst
    umax_877 <= shr_714 when (tmp80_720(0) /=  '0') else type_cast_875_wire_constant;
    addr_of_749_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_749_final_reg_req_0;
      addr_of_749_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_749_final_reg_req_1;
      addr_of_749_final_reg_ack_1<= rack(0);
      addr_of_749_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_749_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_748_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_750,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_932_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_932_final_reg_req_0;
      addr_of_932_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_932_final_reg_req_1;
      addr_of_932_final_reg_ack_1<= rack(0);
      addr_of_932_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_932_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_931_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidxx_xi_933,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    array_obj_ref_1128_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= array_obj_ref_1128_final_reg_req_0;
      array_obj_ref_1128_final_reg_ack_0<= wack(0);
      rreq(0) <= array_obj_ref_1128_final_reg_req_1;
      array_obj_ref_1128_final_reg_ack_1<= rack(0);
      array_obj_ref_1128_final_reg : InterlockBuffer generic map ( -- 
        name => "array_obj_ref_1128_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1128_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx43x_xi_1129,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    array_obj_ref_1140_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= array_obj_ref_1140_final_reg_req_0;
      array_obj_ref_1140_final_reg_ack_0<= wack(0);
      rreq(0) <= array_obj_ref_1140_final_reg_req_1;
      array_obj_ref_1140_final_reg_ack_1<= rack(0);
      array_obj_ref_1140_final_reg : InterlockBuffer generic map ( -- 
        name => "array_obj_ref_1140_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1140_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx48x_xi_1141,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1009_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1009_inst_req_0;
      type_cast_1009_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1009_inst_req_1;
      type_cast_1009_inst_ack_1<= rack(0);
      type_cast_1009_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1009_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr19x_xi_1006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22x_xi_1010,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1030_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1030_inst_req_0;
      type_cast_1030_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1030_inst_req_1;
      type_cast_1030_inst_ack_1<= rack(0);
      type_cast_1030_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1030_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr25x_xi_1027,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28x_xi_1031,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1051_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1051_inst_req_0;
      type_cast_1051_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1051_inst_req_1;
      type_cast_1051_inst_ack_1<= rack(0);
      type_cast_1051_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1051_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr31x_xi_1048,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34x_xi_1052,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1116_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1116_inst_req_0;
      type_cast_1116_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1116_inst_req_1;
      type_cast_1116_inst_ack_1<= rack(0);
      type_cast_1116_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1116_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnextx_xi_1161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1116_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_742_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_742_inst_req_0;
      type_cast_742_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_742_inst_req_1;
      type_cast_742_inst_ack_1<= rack(0);
      type_cast_742_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_742_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_858,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_742_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_757_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_757_inst_req_0;
      type_cast_757_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_757_inst_req_1;
      type_cast_757_inst_ack_1<= rack(0);
      type_cast_757_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_757_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_754,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_758,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_767_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_767_inst_req_0;
      type_cast_767_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_767_inst_req_1;
      type_cast_767_inst_ack_1<= rack(0);
      type_cast_767_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_767_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr11_764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv14_768,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_777_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_777_inst_req_0;
      type_cast_777_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_777_inst_req_1;
      type_cast_777_inst_ack_1<= rack(0);
      type_cast_777_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_777_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr17_774,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_778,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_787_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_787_inst_req_0;
      type_cast_787_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_787_inst_req_1;
      type_cast_787_inst_ack_1<= rack(0);
      type_cast_787_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_787_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr23_784,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_788,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_797_inst_req_0;
      type_cast_797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_797_inst_req_1;
      type_cast_797_inst_ack_1<= rack(0);
      type_cast_797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr29_794,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_798,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_807_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_807_inst_req_0;
      type_cast_807_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_807_inst_req_1;
      type_cast_807_inst_ack_1<= rack(0);
      type_cast_807_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_807_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr35_804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_808,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_817_inst_req_0;
      type_cast_817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_817_inst_req_1;
      type_cast_817_inst_ack_1<= rack(0);
      type_cast_817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr41_814,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_827_inst_req_0;
      type_cast_827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_827_inst_req_1;
      type_cast_827_inst_ack_1<= rack(0);
      type_cast_827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_827_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr47_824,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_828,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_887_inst
    process(tmp81_883) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp81_883(63 downto 0);
      type_cast_887_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_892_inst
    process(ASHR_i64_i64_891_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_891_wire(63 downto 0);
      phitmp_893 <= tmp_var; -- 
    end process;
    type_cast_899_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_899_inst_req_0;
      type_cast_899_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_899_inst_req_1;
      type_cast_899_inst_ack_1<= rack(0);
      type_cast_899_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_899_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_893,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_899_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_925_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_925_inst_req_0;
      type_cast_925_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_925_inst_req_1;
      type_cast_925_inst_ack_1<= rack(0);
      type_cast_925_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_925_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => and70_909,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_926,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_946_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_946_inst_req_0;
      type_cast_946_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_946_inst_req_1;
      type_cast_946_inst_ack_1<= rack(0);
      type_cast_946_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_946_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xi_943,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_947,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_967_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_967_inst_req_0;
      type_cast_967_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_967_inst_req_1;
      type_cast_967_inst_ack_1<= rack(0);
      type_cast_967_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_967_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr7x_xi_964,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10x_xi_968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_988_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_988_inst_req_0;
      type_cast_988_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_988_inst_req_1;
      type_cast_988_inst_ack_1<= rack(0);
      type_cast_988_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_988_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr13x_xi_985,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16x_xi_989,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1128_index_1_rename
    process(R_tmp2_1127_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp2_1127_resized;
      ov(2 downto 0) := iv;
      R_tmp2_1127_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1128_index_1_resize
    process(tmp2_1123) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp2_1123;
      ov := iv(2 downto 0);
      R_tmp2_1127_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1128_root_address_inst
    process(array_obj_ref_1128_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1128_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_1128_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1140_index_1_rename
    process(R_tmp3_1139_resized) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_tmp3_1139_resized;
      ov(2 downto 0) := iv;
      R_tmp3_1139_scaled <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1140_index_1_resize
    process(tmp3_1135) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp3_1135;
      ov := iv(2 downto 0);
      R_tmp3_1139_resized <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1140_root_address_inst
    process(array_obj_ref_1140_final_offset) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1140_final_offset;
      ov(2 downto 0) := iv;
      array_obj_ref_1140_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_748_index_1_rename
    process(R_indvar_747_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_747_resized;
      ov(13 downto 0) := iv;
      R_indvar_747_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_748_index_1_resize
    process(indvar_736) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_736;
      ov := iv(13 downto 0);
      R_indvar_747_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_748_root_address_inst
    process(array_obj_ref_748_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_748_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_748_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_931_index_1_rename
    process(R_ix_x0x_xlcssa_930_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_930_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_930_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_931_index_1_resize
    process(ix_x0x_xlcssa_896) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_896;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_930_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_931_root_address_inst
    process(array_obj_ref_931_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_931_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_931_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1019_addr_0
    process(ptr_deref_1019_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1019_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1019_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1019_base_resize
    process(arrayidx23x_xi_1017) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx23x_xi_1017;
      ov := iv(2 downto 0);
      ptr_deref_1019_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1019_gather_scatter
    process(conv22x_xi_1010) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv22x_xi_1010;
      ov(7 downto 0) := iv;
      ptr_deref_1019_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1019_root_address_inst
    process(ptr_deref_1019_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1019_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1019_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1040_addr_0
    process(ptr_deref_1040_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1040_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1040_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1040_base_resize
    process(arrayidx29x_xi_1038) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx29x_xi_1038;
      ov := iv(2 downto 0);
      ptr_deref_1040_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1040_gather_scatter
    process(conv28x_xi_1031) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv28x_xi_1031;
      ov(7 downto 0) := iv;
      ptr_deref_1040_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1040_root_address_inst
    process(ptr_deref_1040_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1040_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1040_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1061_addr_0
    process(ptr_deref_1061_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1061_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1061_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1061_base_resize
    process(arrayidx35x_xi_1059) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx35x_xi_1059;
      ov := iv(2 downto 0);
      ptr_deref_1061_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1061_gather_scatter
    process(conv34x_xi_1052) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv34x_xi_1052;
      ov(7 downto 0) := iv;
      ptr_deref_1061_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1061_root_address_inst
    process(ptr_deref_1061_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1061_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1061_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1144_addr_0
    process(ptr_deref_1144_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1144_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1144_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1144_base_resize
    process(arrayidx43x_xi_1129) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx43x_xi_1129;
      ov := iv(2 downto 0);
      ptr_deref_1144_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1144_gather_scatter
    process(ptr_deref_1144_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1144_data_0;
      ov(7 downto 0) := iv;
      tmp44x_xi_1145 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1144_root_address_inst
    process(ptr_deref_1144_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1144_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1144_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1151_addr_0
    process(ptr_deref_1151_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1151_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_1151_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1151_base_resize
    process(arrayidx48x_xi_1141) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx48x_xi_1141;
      ov := iv(2 downto 0);
      ptr_deref_1151_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1151_gather_scatter
    process(ptr_deref_1151_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1151_data_0;
      ov(7 downto 0) := iv;
      tmp49x_xi_1152 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1151_root_address_inst
    process(ptr_deref_1151_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1151_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_1151_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_753_addr_0
    process(ptr_deref_753_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_753_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_753_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_753_base_resize
    process(arrayidx_750) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_750;
      ov := iv(13 downto 0);
      ptr_deref_753_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_753_gather_scatter
    process(ptr_deref_753_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_753_data_0;
      ov(63 downto 0) := iv;
      tmp5_754 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_753_root_address_inst
    process(ptr_deref_753_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_753_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_753_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_addr_0
    process(ptr_deref_936_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_936_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_base_resize
    process(arrayidxx_xi_933) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidxx_xi_933;
      ov := iv(13 downto 0);
      ptr_deref_936_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_gather_scatter
    process(ptr_deref_936_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_data_0;
      ov(63 downto 0) := iv;
      tmp1x_xi_937 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_936_root_address_inst
    process(ptr_deref_936_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_936_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_936_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_956_addr_0
    process(ptr_deref_956_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_956_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_956_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_956_base_resize
    process(arrayidx5x_xi_954) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx5x_xi_954;
      ov := iv(2 downto 0);
      ptr_deref_956_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_956_gather_scatter
    process(convx_xi_947) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := convx_xi_947;
      ov(7 downto 0) := iv;
      ptr_deref_956_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_956_root_address_inst
    process(ptr_deref_956_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_956_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_956_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_977_addr_0
    process(ptr_deref_977_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_977_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_977_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_977_base_resize
    process(arrayidx11x_xi_975) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx11x_xi_975;
      ov := iv(2 downto 0);
      ptr_deref_977_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_977_gather_scatter
    process(conv10x_xi_968) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv10x_xi_968;
      ov(7 downto 0) := iv;
      ptr_deref_977_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_977_root_address_inst
    process(ptr_deref_977_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_977_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_977_root_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_998_addr_0
    process(ptr_deref_998_root_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_998_root_address;
      ov(2 downto 0) := iv;
      ptr_deref_998_word_address_0 <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_998_base_resize
    process(arrayidx17x_xi_996) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx17x_xi_996;
      ov := iv(2 downto 0);
      ptr_deref_998_resized_base_address <= ov(2 downto 0);
      --
    end process;
    -- equivalence ptr_deref_998_gather_scatter
    process(conv16x_xi_989) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv16x_xi_989;
      ov(7 downto 0) := iv;
      ptr_deref_998_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_998_root_address_inst
    process(ptr_deref_998_resized_base_address) --
      variable iv : std_logic_vector(2 downto 0);
      variable ov : std_logic_vector(2 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_998_resized_base_address;
      ov(2 downto 0) := iv;
      ptr_deref_998_root_address <= ov(2 downto 0);
      --
    end process;
    if_stmt_1070_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp53x_xi_1069;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1070_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1070_branch_req_0,
          ack0 => if_stmt_1070_branch_ack_0,
          ack1 => if_stmt_1070_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1167_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1166;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1167_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1167_branch_req_0,
          ack0 => if_stmt_1167_branch_ack_0,
          ack1 => if_stmt_1167_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_702_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_701;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_702_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_702_branch_req_0,
          ack0 => if_stmt_702_branch_ack_0,
          ack1 => if_stmt_702_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_864_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_863;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_864_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_864_branch_req_0,
          ack0 => if_stmt_864_branch_ack_0,
          ack1 => if_stmt_864_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_916_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_915;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_916_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_916_branch_req_0,
          ack0 => if_stmt_916_branch_ack_0,
          ack1 => if_stmt_916_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1087_inst
    process(and70_909) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(and70_909, type_cast_1086_wire_constant, tmp_var);
      tmpx_xopx_xi_1088 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1099_inst
    process(iNsTr_29_1094) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_29_1094, type_cast_1098_wire_constant, tmp_var);
      xx_xopx_xi_1100 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1134_inst
    process(tmp2_1123) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_1123, type_cast_1133_wire_constant, tmp_var);
      tmp3_1135 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1160_inst
    process(indvarx_xi_1110) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvarx_xi_1110, type_cast_1159_wire_constant, tmp_var);
      indvarx_xnextx_xi_1161 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_857_inst
    process(indvar_736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_736, type_cast_856_wire_constant, tmp_var);
      indvarx_xnext_858 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1093_inst
    process(tmpx_xopx_xi_1088) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tmpx_xopx_xi_1088, type_cast_1092_wire_constant, tmp_var);
      iNsTr_29_1094 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_908_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(size_buffer, type_cast_907_wire_constant, tmp_var);
      and70_909 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_891_inst
    process(type_cast_887_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_887_wire, type_cast_890_wire_constant, tmp_var);
      ASHR_i64_i64_891_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1068_inst
    process(conv74_926) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv74_926, type_cast_1067_wire_constant, tmp_var);
      cmp53x_xi_1069 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1165_inst
    process(indvarx_xnextx_xi_1161, tmp58x_xi_1107) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnextx_xi_1161, tmp58x_xi_1107, tmp_var);
      exitcond1_1166 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_862_inst
    process(indvarx_xnext_858, umax4_733) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_858, umax4_733, tmp_var);
      exitcond_863 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_914_inst
    process(and70_909) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and70_909, type_cast_913_wire_constant, tmp_var);
      tobool_915 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1005_inst
    process(tmp1x_xi_937) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_937, type_cast_1004_wire_constant, tmp_var);
      shr19x_xi_1006 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1026_inst
    process(tmp1x_xi_937) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_937, type_cast_1025_wire_constant, tmp_var);
      shr25x_xi_1027 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1047_inst
    process(tmp1x_xi_937) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_937, type_cast_1046_wire_constant, tmp_var);
      shr31x_xi_1048 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_713_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_712_wire_constant, tmp_var);
      shr_714 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_763_inst
    process(tmp5_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_754, type_cast_762_wire_constant, tmp_var);
      shr11_764 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_773_inst
    process(tmp5_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_754, type_cast_772_wire_constant, tmp_var);
      shr17_774 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_783_inst
    process(tmp5_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_754, type_cast_782_wire_constant, tmp_var);
      shr23_784 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_793_inst
    process(tmp5_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_754, type_cast_792_wire_constant, tmp_var);
      shr29_794 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_803_inst
    process(tmp5_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_754, type_cast_802_wire_constant, tmp_var);
      shr35_804 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_813_inst
    process(tmp5_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_754, type_cast_812_wire_constant, tmp_var);
      shr41_814 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_823_inst
    process(tmp5_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp5_754, type_cast_822_wire_constant, tmp_var);
      shr47_824 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_942_inst
    process(tmp1x_xi_937) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_937, type_cast_941_wire_constant, tmp_var);
      shrx_xi_943 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_963_inst
    process(tmp1x_xi_937) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_937, type_cast_962_wire_constant, tmp_var);
      shr7x_xi_964 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_984_inst
    process(tmp1x_xi_937) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1x_xi_937, type_cast_983_wire_constant, tmp_var);
      shr13x_xi_985 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1122_inst
    process(indvarx_xi_1110) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvarx_xi_1110, type_cast_1121_wire_constant, tmp_var);
      tmp2_1123 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_882_inst
    process(umax_877) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_877, type_cast_881_wire_constant, tmp_var);
      tmp81_883 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_1081_inst
    process(conv74_926) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv74_926, type_cast_1080_wire_constant, tmp_var);
      tmp55x_xi_1082 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_700_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_699_wire_constant, tmp_var);
      cmp77_701 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_719_inst
    process(shr_714) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_714, type_cast_718_wire_constant, tmp_var);
      tmp80_720 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_725_inst
    process(shr_714) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_714, type_cast_724_wire_constant, tmp_var);
      tmp_726 <= tmp_var; --
    end process;
    -- shared split operator group (32) : array_obj_ref_1128_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_tmp2_1127_scaled;
      array_obj_ref_1128_final_offset <= data_out(2 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1128_index_offset_req_0;
      array_obj_ref_1128_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1128_index_offset_req_1;
      array_obj_ref_1128_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : array_obj_ref_1140_index_offset 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(2 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_tmp3_1139_scaled;
      array_obj_ref_1140_final_offset <= data_out(2 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1140_index_offset_req_0;
      array_obj_ref_1140_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1140_index_offset_req_1;
      array_obj_ref_1140_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 3,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : array_obj_ref_748_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_747_scaled;
      array_obj_ref_748_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_748_index_offset_req_0;
      array_obj_ref_748_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_748_index_offset_req_1;
      array_obj_ref_748_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_931_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_930_scaled;
      array_obj_ref_931_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_931_index_offset_req_0;
      array_obj_ref_931_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_931_index_offset_req_1;
      array_obj_ref_931_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared load operator group (0) : ptr_deref_1144_load_0 ptr_deref_1151_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1144_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1151_load_0_req_0;
      ptr_deref_1144_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1151_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1144_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1151_load_0_req_1;
      ptr_deref_1144_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1151_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1144_word_address_0 & ptr_deref_1151_word_address_0;
      ptr_deref_1144_data_0 <= data_out(15 downto 8);
      ptr_deref_1151_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 3,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(2 downto 0),
          mtag => memory_space_3_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_936_load_0 ptr_deref_753_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_936_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_753_load_0_req_0;
      ptr_deref_936_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_753_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_936_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_753_load_0_req_1;
      ptr_deref_936_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_753_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_936_word_address_0 & ptr_deref_753_word_address_0;
      ptr_deref_936_data_0 <= data_out(127 downto 64);
      ptr_deref_753_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : ptr_deref_998_store_0 ptr_deref_1019_store_0 ptr_deref_977_store_0 ptr_deref_956_store_0 ptr_deref_1040_store_0 ptr_deref_1061_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(17 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_998_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1019_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_977_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_956_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1040_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1061_store_0_req_0;
      ptr_deref_998_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1019_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_977_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_956_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1040_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1061_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_998_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1019_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_977_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_956_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1040_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1061_store_0_req_1;
      ptr_deref_998_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1019_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_977_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_956_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1040_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1061_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_998_word_address_0 & ptr_deref_1019_word_address_0 & ptr_deref_977_word_address_0 & ptr_deref_956_word_address_0 & ptr_deref_1040_word_address_0 & ptr_deref_1061_word_address_0;
      data_in <= ptr_deref_998_data_0 & ptr_deref_1019_data_0 & ptr_deref_977_data_0 & ptr_deref_956_data_0 & ptr_deref_1040_data_0 & ptr_deref_1061_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 3,
        data_width => 8,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(2 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 6,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_829_inst WPIPE_maxpool_output_pipe_832_inst WPIPE_maxpool_output_pipe_835_inst WPIPE_maxpool_output_pipe_838_inst WPIPE_maxpool_output_pipe_850_inst WPIPE_maxpool_output_pipe_847_inst WPIPE_maxpool_output_pipe_1146_inst WPIPE_maxpool_output_pipe_1153_inst WPIPE_maxpool_output_pipe_844_inst WPIPE_maxpool_output_pipe_841_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal sample_req, sample_ack : BooleanArray( 9 downto 0);
      signal update_req, update_ack : BooleanArray( 9 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 9 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_829_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_832_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_835_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_838_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_850_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_847_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1146_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1153_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_844_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_841_inst_req_0;
      WPIPE_maxpool_output_pipe_829_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_832_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_835_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_838_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_850_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_847_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1146_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1153_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_844_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_841_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_829_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_832_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_835_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_838_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_850_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_847_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1146_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1153_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_844_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_841_inst_req_1;
      WPIPE_maxpool_output_pipe_829_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_832_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_835_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_838_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_850_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_847_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1146_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1153_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_844_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_841_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      data_in <= conv50_828 & conv44_818 & conv38_808 & conv32_798 & conv8_758 & conv14_768 & tmp44x_xi_1145 & tmp49x_xi_1152 & conv20_778 & conv26_788;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 10, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 1,
      addr_width => 3,
      data_width => 8,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 3,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendModule is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
    output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendModule;
architecture sendModule_arch of sendModule is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendModule_CP_7961_start: Boolean;
  signal sendModule_CP_7961_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_3214_req_0 : boolean;
  signal type_cast_3280_inst_ack_1 : boolean;
  signal ptr_deref_3339_load_0_req_1 : boolean;
  signal ptr_deref_3339_load_0_ack_1 : boolean;
  signal ptr_deref_3335_load_0_req_0 : boolean;
  signal phi_stmt_3214_ack_0 : boolean;
  signal ptr_deref_3335_load_0_ack_0 : boolean;
  signal array_obj_ref_3330_index_offset_req_1 : boolean;
  signal array_obj_ref_3330_index_offset_ack_1 : boolean;
  signal SUB_u16_u16_3233_inst_req_0 : boolean;
  signal SUB_u16_u16_3233_inst_ack_0 : boolean;
  signal ptr_deref_3335_load_0_req_1 : boolean;
  signal n_col_3249_3218_buf_req_0 : boolean;
  signal n_col_3249_3218_buf_ack_0 : boolean;
  signal array_obj_ref_3330_index_offset_ack_0 : boolean;
  signal ptr_deref_3339_load_0_req_0 : boolean;
  signal ptr_deref_3339_load_0_ack_0 : boolean;
  signal RPIPE_output_pipe_3342_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3342_inst_ack_1 : boolean;
  signal RPIPE_output_pipe_3342_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3342_inst_ack_0 : boolean;
  signal type_cast_3271_inst_ack_1 : boolean;
  signal phi_stmt_3214_req_1 : boolean;
  signal type_cast_3271_inst_req_1 : boolean;
  signal array_obj_ref_3330_index_offset_req_0 : boolean;
  signal ptr_deref_3335_load_0_ack_1 : boolean;
  signal array_obj_ref_3320_index_offset_ack_1 : boolean;
  signal type_cast_3271_inst_ack_0 : boolean;
  signal type_cast_3271_inst_req_0 : boolean;
  signal type_cast_3280_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3183_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3183_inst_ack_0 : boolean;
  signal addr_of_3331_final_reg_ack_1 : boolean;
  signal RPIPE_output_pipe_3183_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3183_inst_ack_1 : boolean;
  signal n_row_3260_3223_buf_ack_1 : boolean;
  signal addr_of_3331_final_reg_req_1 : boolean;
  signal RPIPE_output_pipe_3186_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3186_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3186_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3186_inst_ack_1 : boolean;
  signal n_row_3260_3223_buf_req_1 : boolean;
  signal type_cast_3280_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3189_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3189_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3189_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3189_inst_ack_1 : boolean;
  signal do_while_stmt_3197_branch_req_0 : boolean;
  signal array_obj_ref_3320_index_offset_req_1 : boolean;
  signal n_row_3260_3223_buf_ack_0 : boolean;
  signal SUB_u16_u16_3233_inst_ack_1 : boolean;
  signal array_obj_ref_3320_index_offset_ack_0 : boolean;
  signal n_row_3260_3223_buf_req_0 : boolean;
  signal addr_of_3321_final_reg_ack_1 : boolean;
  signal type_cast_3280_inst_req_0 : boolean;
  signal phi_stmt_3199_req_1 : boolean;
  signal addr_of_3321_final_reg_req_1 : boolean;
  signal phi_stmt_3199_req_0 : boolean;
  signal addr_of_3321_final_reg_ack_0 : boolean;
  signal addr_of_3331_final_reg_ack_0 : boolean;
  signal array_obj_ref_3320_index_offset_req_0 : boolean;
  signal phi_stmt_3199_ack_0 : boolean;
  signal addr_of_3321_final_reg_req_0 : boolean;
  signal phi_stmt_3219_ack_0 : boolean;
  signal n_chl_3268_3213_buf_ack_1 : boolean;
  signal phi_stmt_3219_req_0 : boolean;
  signal phi_stmt_3219_req_1 : boolean;
  signal addr_of_3331_final_reg_req_0 : boolean;
  signal n_address1_3298_3203_buf_req_0 : boolean;
  signal SUB_u16_u16_3233_inst_req_1 : boolean;
  signal n_address1_3298_3203_buf_ack_0 : boolean;
  signal n_address1_3298_3203_buf_req_1 : boolean;
  signal n_address1_3298_3203_buf_ack_1 : boolean;
  signal n_col_3249_3218_buf_ack_1 : boolean;
  signal n_col_3249_3218_buf_req_1 : boolean;
  signal ptr_deref_3516_store_0_req_0 : boolean;
  signal phi_stmt_3204_req_1 : boolean;
  signal phi_stmt_3204_req_0 : boolean;
  signal ptr_deref_3516_store_0_ack_0 : boolean;
  signal phi_stmt_3204_ack_0 : boolean;
  signal type_cast_3207_inst_req_0 : boolean;
  signal type_cast_3207_inst_ack_0 : boolean;
  signal type_cast_3207_inst_req_1 : boolean;
  signal type_cast_3207_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3540_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3540_inst_ack_0 : boolean;
  signal n_address2_3312_3208_buf_req_0 : boolean;
  signal n_address2_3312_3208_buf_ack_0 : boolean;
  signal n_address2_3312_3208_buf_req_1 : boolean;
  signal n_address2_3312_3208_buf_ack_1 : boolean;
  signal phi_stmt_3209_req_1 : boolean;
  signal phi_stmt_3209_req_0 : boolean;
  signal phi_stmt_3209_ack_0 : boolean;
  signal n_chl_3268_3213_buf_req_0 : boolean;
  signal n_chl_3268_3213_buf_ack_0 : boolean;
  signal n_chl_3268_3213_buf_req_1 : boolean;
  signal RPIPE_output_pipe_3345_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3345_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3345_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3345_inst_ack_1 : boolean;
  signal slice_3349_inst_req_0 : boolean;
  signal slice_3349_inst_ack_0 : boolean;
  signal slice_3349_inst_req_1 : boolean;
  signal slice_3349_inst_ack_1 : boolean;
  signal slice_3353_inst_req_0 : boolean;
  signal slice_3353_inst_ack_0 : boolean;
  signal slice_3353_inst_req_1 : boolean;
  signal slice_3353_inst_ack_1 : boolean;
  signal slice_3357_inst_req_0 : boolean;
  signal slice_3357_inst_ack_0 : boolean;
  signal slice_3357_inst_req_1 : boolean;
  signal slice_3357_inst_ack_1 : boolean;
  signal ptr_deref_3516_store_0_ack_1 : boolean;
  signal slice_3361_inst_req_0 : boolean;
  signal slice_3361_inst_ack_0 : boolean;
  signal slice_3361_inst_req_1 : boolean;
  signal slice_3361_inst_ack_1 : boolean;
  signal slice_3365_inst_req_0 : boolean;
  signal slice_3365_inst_ack_0 : boolean;
  signal slice_3365_inst_req_1 : boolean;
  signal slice_3365_inst_ack_1 : boolean;
  signal slice_3369_inst_req_0 : boolean;
  signal slice_3369_inst_ack_0 : boolean;
  signal slice_3369_inst_req_1 : boolean;
  signal slice_3369_inst_ack_1 : boolean;
  signal do_while_stmt_3197_branch_ack_1 : boolean;
  signal slice_3373_inst_req_0 : boolean;
  signal slice_3373_inst_ack_0 : boolean;
  signal slice_3373_inst_req_1 : boolean;
  signal slice_3373_inst_ack_1 : boolean;
  signal slice_3377_inst_req_0 : boolean;
  signal slice_3377_inst_ack_0 : boolean;
  signal slice_3377_inst_req_1 : boolean;
  signal slice_3377_inst_ack_1 : boolean;
  signal do_while_stmt_3197_branch_ack_0 : boolean;
  signal ptr_deref_3516_store_0_req_1 : boolean;
  signal EQ_u2_u1_3390_inst_req_0 : boolean;
  signal EQ_u2_u1_3390_inst_ack_0 : boolean;
  signal EQ_u2_u1_3390_inst_req_1 : boolean;
  signal EQ_u2_u1_3390_inst_ack_1 : boolean;
  signal W_output_data1_3262_delayed_14_0_3392_inst_req_0 : boolean;
  signal W_output_data1_3262_delayed_14_0_3392_inst_ack_0 : boolean;
  signal W_output_data1_3262_delayed_14_0_3392_inst_req_1 : boolean;
  signal W_output_data1_3262_delayed_14_0_3392_inst_ack_1 : boolean;
  signal EQ_u2_u1_3404_inst_req_0 : boolean;
  signal EQ_u2_u1_3404_inst_ack_0 : boolean;
  signal EQ_u2_u1_3404_inst_req_1 : boolean;
  signal EQ_u2_u1_3404_inst_ack_1 : boolean;
  signal SUB_u16_u16_3528_inst_ack_1 : boolean;
  signal W_output_data1_3270_delayed_14_0_3406_inst_req_0 : boolean;
  signal W_output_data1_3270_delayed_14_0_3406_inst_ack_0 : boolean;
  signal W_output_data1_3270_delayed_14_0_3406_inst_req_1 : boolean;
  signal W_output_data1_3270_delayed_14_0_3406_inst_ack_1 : boolean;
  signal SUB_u16_u16_3528_inst_req_1 : boolean;
  signal EQ_u2_u1_3418_inst_req_0 : boolean;
  signal EQ_u2_u1_3418_inst_ack_0 : boolean;
  signal EQ_u2_u1_3418_inst_req_1 : boolean;
  signal EQ_u2_u1_3418_inst_ack_1 : boolean;
  signal SUB_u16_u16_3528_inst_ack_0 : boolean;
  signal W_output_data1_3278_delayed_14_0_3420_inst_req_0 : boolean;
  signal W_output_data1_3278_delayed_14_0_3420_inst_ack_0 : boolean;
  signal W_output_data1_3278_delayed_14_0_3420_inst_req_1 : boolean;
  signal W_output_data1_3278_delayed_14_0_3420_inst_ack_1 : boolean;
  signal SUB_u16_u16_3528_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3540_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3540_inst_req_1 : boolean;
  signal EQ_u2_u1_3432_inst_req_0 : boolean;
  signal EQ_u2_u1_3432_inst_ack_0 : boolean;
  signal EQ_u2_u1_3432_inst_req_1 : boolean;
  signal EQ_u2_u1_3432_inst_ack_1 : boolean;
  signal W_output_data1_3286_delayed_14_0_3434_inst_req_0 : boolean;
  signal W_output_data1_3286_delayed_14_0_3434_inst_ack_0 : boolean;
  signal W_output_data1_3286_delayed_14_0_3434_inst_req_1 : boolean;
  signal W_output_data1_3286_delayed_14_0_3434_inst_ack_1 : boolean;
  signal EQ_u2_u1_3446_inst_req_0 : boolean;
  signal EQ_u2_u1_3446_inst_ack_0 : boolean;
  signal EQ_u2_u1_3446_inst_req_1 : boolean;
  signal EQ_u2_u1_3446_inst_ack_1 : boolean;
  signal W_output_data2_3294_delayed_14_0_3448_inst_req_0 : boolean;
  signal W_output_data2_3294_delayed_14_0_3448_inst_ack_0 : boolean;
  signal W_output_data2_3294_delayed_14_0_3448_inst_req_1 : boolean;
  signal W_output_data2_3294_delayed_14_0_3448_inst_ack_1 : boolean;
  signal EQ_u2_u1_3460_inst_req_0 : boolean;
  signal EQ_u2_u1_3460_inst_ack_0 : boolean;
  signal EQ_u2_u1_3460_inst_req_1 : boolean;
  signal EQ_u2_u1_3460_inst_ack_1 : boolean;
  signal W_output_data2_3302_delayed_14_0_3462_inst_req_0 : boolean;
  signal W_output_data2_3302_delayed_14_0_3462_inst_ack_0 : boolean;
  signal W_output_data2_3302_delayed_14_0_3462_inst_req_1 : boolean;
  signal W_output_data2_3302_delayed_14_0_3462_inst_ack_1 : boolean;
  signal EQ_u2_u1_3474_inst_req_0 : boolean;
  signal EQ_u2_u1_3474_inst_ack_0 : boolean;
  signal EQ_u2_u1_3474_inst_req_1 : boolean;
  signal EQ_u2_u1_3474_inst_ack_1 : boolean;
  signal W_output_data2_3310_delayed_14_0_3476_inst_req_0 : boolean;
  signal W_output_data2_3310_delayed_14_0_3476_inst_ack_0 : boolean;
  signal W_output_data2_3310_delayed_14_0_3476_inst_req_1 : boolean;
  signal W_output_data2_3310_delayed_14_0_3476_inst_ack_1 : boolean;
  signal EQ_u2_u1_3488_inst_req_0 : boolean;
  signal EQ_u2_u1_3488_inst_ack_0 : boolean;
  signal EQ_u2_u1_3488_inst_req_1 : boolean;
  signal EQ_u2_u1_3488_inst_ack_1 : boolean;
  signal W_output_data2_3318_delayed_14_0_3490_inst_req_0 : boolean;
  signal W_output_data2_3318_delayed_14_0_3490_inst_ack_0 : boolean;
  signal W_output_data2_3318_delayed_14_0_3490_inst_req_1 : boolean;
  signal W_output_data2_3318_delayed_14_0_3490_inst_ack_1 : boolean;
  signal W_fetch_addr1_3322_delayed_8_0_3499_inst_req_0 : boolean;
  signal W_fetch_addr1_3322_delayed_8_0_3499_inst_ack_0 : boolean;
  signal W_fetch_addr1_3322_delayed_8_0_3499_inst_req_1 : boolean;
  signal W_fetch_addr1_3322_delayed_8_0_3499_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3510_inst_req_0 : boolean;
  signal CONCAT_u32_u64_3510_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_3510_inst_req_1 : boolean;
  signal CONCAT_u32_u64_3510_inst_ack_1 : boolean;
  signal ptr_deref_3503_store_0_req_0 : boolean;
  signal ptr_deref_3503_store_0_ack_0 : boolean;
  signal ptr_deref_3503_store_0_req_1 : boolean;
  signal ptr_deref_3503_store_0_ack_1 : boolean;
  signal W_fetch_addr2_3332_delayed_8_0_3512_inst_req_0 : boolean;
  signal W_fetch_addr2_3332_delayed_8_0_3512_inst_ack_0 : boolean;
  signal W_fetch_addr2_3332_delayed_8_0_3512_inst_req_1 : boolean;
  signal W_fetch_addr2_3332_delayed_8_0_3512_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3523_inst_req_0 : boolean;
  signal CONCAT_u32_u64_3523_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_3523_inst_req_1 : boolean;
  signal CONCAT_u32_u64_3523_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendModule_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendModule_CP_7961_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendModule_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_7961_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendModule_CP_7961_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_7961_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendModule_CP_7961: Block -- control-path 
    signal sendModule_CP_7961_elements: BooleanArray(291 downto 0);
    -- 
  begin -- 
    sendModule_CP_7961_elements(0) <= sendModule_CP_7961_start;
    sendModule_CP_7961_symbol <= sendModule_CP_7961_elements(291);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3181/$entry
      -- CP-element group 0: 	 branch_block_stmt_3181/branch_block_stmt_3181__entry__
      -- CP-element group 0: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196__entry__
      -- CP-element group 0: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/$entry
      -- CP-element group 0: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_Sample/rr
      -- 
    rr_7985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(0), ack => RPIPE_output_pipe_3183_inst_req_0); -- 
    -- CP-element group 1:  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	289 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	290 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_3181/do_while_stmt_3197__exit__
      -- CP-element group 1: 	 branch_block_stmt_3181/assign_stmt_3542__entry__
      -- CP-element group 1: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_Sample/req
      -- CP-element group 1: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_3181/assign_stmt_3542/$entry
      -- 
    req_9062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(1), ack => WPIPE_input_done_pipe_3540_inst_req_0); -- 
    sendModule_CP_7961_elements(1) <= sendModule_CP_7961_elements(289);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_update_start_
      -- CP-element group 2: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_Update/cr
      -- 
    ra_7986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3183_inst_ack_0, ack => sendModule_CP_7961_elements(2)); -- 
    cr_7990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(2), ack => RPIPE_output_pipe_3183_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3183_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_Sample/rr
      -- 
    ca_7991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3183_inst_ack_1, ack => sendModule_CP_7961_elements(3)); -- 
    rr_7999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(3), ack => RPIPE_output_pipe_3186_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_update_start_
      -- CP-element group 4: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_Update/cr
      -- 
    ra_8000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3186_inst_ack_0, ack => sendModule_CP_7961_elements(4)); -- 
    cr_8004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(4), ack => RPIPE_output_pipe_3186_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3186_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_Sample/rr
      -- 
    ca_8005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3186_inst_ack_1, ack => sendModule_CP_7961_elements(5)); -- 
    rr_8013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(5), ack => RPIPE_output_pipe_3189_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_update_start_
      -- CP-element group 6: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_Update/cr
      -- 
    ra_8014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3189_inst_ack_0, ack => sendModule_CP_7961_elements(6)); -- 
    cr_8018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(6), ack => RPIPE_output_pipe_3189_inst_req_1); -- 
    -- CP-element group 7:  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196__exit__
      -- CP-element group 7: 	 branch_block_stmt_3181/do_while_stmt_3197__entry__
      -- CP-element group 7: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/$exit
      -- CP-element group 7: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_3181/assign_stmt_3184_to_assign_stmt_3196/RPIPE_output_pipe_3189_Update/ca
      -- 
    ca_8019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3189_inst_ack_1, ack => sendModule_CP_7961_elements(7)); -- 
    -- CP-element group 8:  transition  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_3181/do_while_stmt_3197/$entry
      -- CP-element group 8: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197__entry__
      -- 
    sendModule_CP_7961_elements(8) <= sendModule_CP_7961_elements(7);
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	289 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197__exit__
      -- 
    -- Element group sendModule_CP_7961_elements(9) is bound as output of CP function.
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3181/do_while_stmt_3197/loop_back
      -- 
    -- Element group sendModule_CP_7961_elements(10) is bound as output of CP function.
    -- CP-element group 11:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	287 
    -- CP-element group 11: 	288 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_3181/do_while_stmt_3197/condition_done
      -- CP-element group 11: 	 branch_block_stmt_3181/do_while_stmt_3197/loop_taken/$entry
      -- CP-element group 11: 	 branch_block_stmt_3181/do_while_stmt_3197/loop_exit/$entry
      -- 
    sendModule_CP_7961_elements(11) <= sendModule_CP_7961_elements(16);
    -- CP-element group 12:  branch  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	286 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_3181/do_while_stmt_3197/loop_body_done
      -- 
    sendModule_CP_7961_elements(12) <= sendModule_CP_7961_elements(286);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	25 
    -- CP-element group 13: 	44 
    -- CP-element group 13: 	65 
    -- CP-element group 13: 	84 
    -- CP-element group 13: 	103 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/back_edge_to_loop_body
      -- 
    sendModule_CP_7961_elements(13) <= sendModule_CP_7961_elements(10);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	27 
    -- CP-element group 14: 	46 
    -- CP-element group 14: 	67 
    -- CP-element group 14: 	86 
    -- CP-element group 14: 	105 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/first_time_through_loop_body
      -- 
    sendModule_CP_7961_elements(14) <= sendModule_CP_7961_elements(8);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	120 
    -- CP-element group 15: 	130 
    -- CP-element group 15: 	136 
    -- CP-element group 15: 	129 
    -- CP-element group 15: 	137 
    -- CP-element group 15: 	116 
    -- CP-element group 15: 	150 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	278 
    -- CP-element group 15: 	282 
    -- CP-element group 15: 	124 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	39 
    -- CP-element group 15: 	59 
    -- CP-element group 15: 	60 
    -- CP-element group 15: 	78 
    -- CP-element group 15: 	79 
    -- CP-element group 15: 	97 
    -- CP-element group 15: 	98 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/$entry
      -- CP-element group 15: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/loop_body_start
      -- 
    -- Element group sendModule_CP_7961_elements(15) is bound as output of CP function.
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	119 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	281 
    -- CP-element group 16: 	282 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/condition_evaluated
      -- 
    condition_evaluated_8034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_8034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(16), ack => do_while_stmt_3197_branch_req_0); -- 
    sendModule_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(119) & sendModule_CP_7961_elements(20) & sendModule_CP_7961_elements(281) & sendModule_CP_7961_elements(282);
      gj_sendModule_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	38 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	78 
    -- CP-element group 17: 	97 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	61 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	99 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/aggregated_phi_sample_req
      -- CP-element group 17: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_sample_start__ps
      -- 
    sendModule_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(21) & sendModule_CP_7961_elements(38) & sendModule_CP_7961_elements(59) & sendModule_CP_7961_elements(78) & sendModule_CP_7961_elements(97) & sendModule_CP_7961_elements(20);
      gj_sendModule_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	23 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	81 
    -- CP-element group 18: 	100 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	121 
    -- CP-element group 18: 	117 
    -- CP-element group 18: 	286 
    -- CP-element group 18: 	125 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	38 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	78 
    -- CP-element group 18: 	97 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/aggregated_phi_sample_ack
      -- CP-element group 18: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_sample_completed_
      -- 
    sendModule_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(23) & sendModule_CP_7961_elements(41) & sendModule_CP_7961_elements(62) & sendModule_CP_7961_elements(81) & sendModule_CP_7961_elements(100);
      gj_sendModule_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	39 
    -- CP-element group 19: 	60 
    -- CP-element group 19: 	79 
    -- CP-element group 19: 	98 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	63 
    -- CP-element group 19: 	82 
    -- CP-element group 19: 	101 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/aggregated_phi_update_req
      -- CP-element group 19: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_update_start__ps
      -- 
    sendModule_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(22) & sendModule_CP_7961_elements(39) & sendModule_CP_7961_elements(60) & sendModule_CP_7961_elements(79) & sendModule_CP_7961_elements(98);
      gj_sendModule_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	64 
    -- CP-element group 20: 	83 
    -- CP-element group 20: 	102 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/aggregated_phi_update_ack
      -- 
    sendModule_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(24) & sendModule_CP_7961_elements(43) & sendModule_CP_7961_elements(64) & sendModule_CP_7961_elements(83) & sendModule_CP_7961_elements(102);
      gj_sendModule_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	119 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	123 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_sample_start_
      -- 
    sendModule_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(119) & sendModule_CP_7961_elements(18) & sendModule_CP_7961_elements(123);
      gj_sendModule_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	131 
    -- CP-element group 22: 	208 
    -- CP-element group 22: 	216 
    -- CP-element group 22: 	200 
    -- CP-element group 22: 	192 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	19 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_update_start_
      -- 
    sendModule_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(131) & sendModule_CP_7961_elements(208) & sendModule_CP_7961_elements(216) & sendModule_CP_7961_elements(200) & sendModule_CP_7961_elements(192);
      gj_sendModule_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	18 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7961_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	131 
    -- CP-element group 24: 	20 
    -- CP-element group 24: 	214 
    -- CP-element group 24: 	198 
    -- CP-element group 24: 	206 
    -- CP-element group 24: 	190 
    -- CP-element group 24:  members (15) 
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_scale_1/scale_rename_req
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_scale_1/scale_rename_ack
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_resized_1
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_scaled_1
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_scale_1/$exit
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_scale_1/$entry
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_resize_1/index_resize_ack
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_resize_1/index_resize_req
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_resize_1/$exit
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_resize_1/$entry
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_index_computed_1
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_Sample/req
      -- CP-element group 24: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_Sample/$entry
      -- 
    req_8336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(24), ack => array_obj_ref_3320_index_offset_req_0); -- 
    -- Element group sendModule_CP_7961_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	13 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_loopback_trigger
      -- 
    sendModule_CP_7961_elements(25) <= sendModule_CP_7961_elements(13);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_loopback_sample_req
      -- CP-element group 26: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_loopback_sample_req_ps
      -- 
    phi_stmt_3199_loopback_sample_req_8049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3199_loopback_sample_req_8049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(26), ack => phi_stmt_3199_req_1); -- 
    -- Element group sendModule_CP_7961_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	14 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_entry_trigger
      -- 
    sendModule_CP_7961_elements(27) <= sendModule_CP_7961_elements(14);
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_entry_sample_req
      -- CP-element group 28: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_entry_sample_req_ps
      -- 
    phi_stmt_3199_entry_sample_req_8052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3199_entry_sample_req_8052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(28), ack => phi_stmt_3199_req_0); -- 
    -- Element group sendModule_CP_7961_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_phi_mux_ack
      -- CP-element group 29: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3199_phi_mux_ack_ps
      -- 
    phi_stmt_3199_phi_mux_ack_8055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3199_ack_0, ack => sendModule_CP_7961_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3202_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3202_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3202_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3202_sample_completed_
      -- 
    -- Element group sendModule_CP_7961_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3202_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3202_update_start_
      -- 
    -- Element group sendModule_CP_7961_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3202_update_completed__ps
      -- 
    sendModule_CP_7961_elements(32) <= sendModule_CP_7961_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3202_update_completed_
      -- 
    -- Element group sendModule_CP_7961_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => sendModule_CP_7961_elements(31), ack => sendModule_CP_7961_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_Sample/req
      -- 
    req_8076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(34), ack => n_address1_3298_3203_buf_req_0); -- 
    -- Element group sendModule_CP_7961_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_update_start_
      -- CP-element group 35: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_Update/req
      -- 
    req_8081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(35), ack => n_address1_3298_3203_buf_req_1); -- 
    -- Element group sendModule_CP_7961_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_Sample/ack
      -- 
    ack_8077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_3298_3203_buf_ack_0, ack => sendModule_CP_7961_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address1_3203_Update/ack
      -- 
    ack_8082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_3298_3203_buf_ack_1, ack => sendModule_CP_7961_elements(37)); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	119 
    -- CP-element group 38: 	127 
    -- CP-element group 38: 	18 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	17 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_sample_start_
      -- 
    sendModule_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(119) & sendModule_CP_7961_elements(127) & sendModule_CP_7961_elements(18);
      gj_sendModule_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	15 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	138 
    -- CP-element group 39: 	240 
    -- CP-element group 39: 	248 
    -- CP-element group 39: 	224 
    -- CP-element group 39: 	232 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	19 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_update_start_
      -- 
    sendModule_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(138) & sendModule_CP_7961_elements(240) & sendModule_CP_7961_elements(248) & sendModule_CP_7961_elements(224) & sendModule_CP_7961_elements(232);
      gj_sendModule_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	17 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_sample_start__ps
      -- 
    sendModule_CP_7961_elements(40) <= sendModule_CP_7961_elements(17);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	18 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7961_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_update_start__ps
      -- 
    sendModule_CP_7961_elements(42) <= sendModule_CP_7961_elements(19);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	138 
    -- CP-element group 43: 	20 
    -- CP-element group 43: 	238 
    -- CP-element group 43: 	246 
    -- CP-element group 43: 	222 
    -- CP-element group 43: 	230 
    -- CP-element group 43:  members (15) 
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_scale_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_Sample/req
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_update_completed__ps
      -- 
    req_8382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(43), ack => array_obj_ref_3330_index_offset_req_0); -- 
    -- Element group sendModule_CP_7961_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	13 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_loopback_trigger
      -- 
    sendModule_CP_7961_elements(44) <= sendModule_CP_7961_elements(13);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_loopback_sample_req_ps
      -- 
    phi_stmt_3204_loopback_sample_req_8093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3204_loopback_sample_req_8093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(45), ack => phi_stmt_3204_req_1); -- 
    -- Element group sendModule_CP_7961_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	14 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_entry_trigger
      -- 
    sendModule_CP_7961_elements(46) <= sendModule_CP_7961_elements(14);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_entry_sample_req
      -- CP-element group 47: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_entry_sample_req_ps
      -- 
    phi_stmt_3204_entry_sample_req_8096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3204_entry_sample_req_8096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(47), ack => phi_stmt_3204_req_0); -- 
    -- Element group sendModule_CP_7961_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_phi_mux_ack
      -- CP-element group 48: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3204_phi_mux_ack_ps
      -- 
    phi_stmt_3204_phi_mux_ack_8099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3204_ack_0, ack => sendModule_CP_7961_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_sample_start__ps
      -- 
    -- Element group sendModule_CP_7961_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_update_start__ps
      -- 
    -- Element group sendModule_CP_7961_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_Sample/rr
      -- 
    rr_8112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(51), ack => type_cast_3207_inst_req_0); -- 
    sendModule_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(49) & sendModule_CP_7961_elements(53);
      gj_sendModule_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_update_start_
      -- CP-element group 52: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_Update/cr
      -- 
    cr_8117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(52), ack => type_cast_3207_inst_req_1); -- 
    sendModule_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(50) & sendModule_CP_7961_elements(54);
      gj_sendModule_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_Sample/ra
      -- 
    ra_8113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3207_inst_ack_0, ack => sendModule_CP_7961_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3207_Update/ca
      -- 
    ca_8118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3207_inst_ack_1, ack => sendModule_CP_7961_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_Sample/req
      -- 
    req_8130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(55), ack => n_address2_3312_3208_buf_req_0); -- 
    -- Element group sendModule_CP_7961_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_update_start__ps
      -- CP-element group 56: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_update_start_
      -- CP-element group 56: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_Update/req
      -- 
    req_8135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(56), ack => n_address2_3312_3208_buf_req_1); -- 
    -- Element group sendModule_CP_7961_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_Sample/ack
      -- 
    ack_8131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_3312_3208_buf_ack_0, ack => sendModule_CP_7961_elements(57)); -- 
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_address2_3208_Update/ack
      -- 
    ack_8136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_3312_3208_buf_ack_1, ack => sendModule_CP_7961_elements(58)); -- 
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	15 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	119 
    -- CP-element group 59: 	18 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_sample_start_
      -- 
    sendModule_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(119) & sendModule_CP_7961_elements(18);
      gj_sendModule_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	15 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	64 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	19 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_update_start_
      -- 
    sendModule_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(64);
      gj_sendModule_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	17 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_sample_start__ps
      -- 
    sendModule_CP_7961_elements(61) <= sendModule_CP_7961_elements(17);
    -- CP-element group 62:  join  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	18 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7961_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_update_start__ps
      -- 
    sendModule_CP_7961_elements(63) <= sendModule_CP_7961_elements(19);
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	20 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	60 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_update_completed__ps
      -- 
    -- Element group sendModule_CP_7961_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	13 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_loopback_trigger
      -- 
    sendModule_CP_7961_elements(65) <= sendModule_CP_7961_elements(13);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_loopback_sample_req
      -- CP-element group 66: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_loopback_sample_req_ps
      -- 
    phi_stmt_3209_loopback_sample_req_8147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3209_loopback_sample_req_8147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(66), ack => phi_stmt_3209_req_1); -- 
    -- Element group sendModule_CP_7961_elements(66) is bound as output of CP function.
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_entry_trigger
      -- 
    sendModule_CP_7961_elements(67) <= sendModule_CP_7961_elements(14);
    -- CP-element group 68:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_entry_sample_req
      -- CP-element group 68: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_entry_sample_req_ps
      -- 
    phi_stmt_3209_entry_sample_req_8150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3209_entry_sample_req_8150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(68), ack => phi_stmt_3209_req_0); -- 
    -- Element group sendModule_CP_7961_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_phi_mux_ack
      -- CP-element group 69: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3209_phi_mux_ack_ps
      -- 
    phi_stmt_3209_phi_mux_ack_8153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3209_ack_0, ack => sendModule_CP_7961_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3212_sample_start__ps
      -- CP-element group 70: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3212_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3212_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3212_sample_completed_
      -- 
    -- Element group sendModule_CP_7961_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3212_update_start__ps
      -- CP-element group 71: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3212_update_start_
      -- 
    -- Element group sendModule_CP_7961_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3212_update_completed__ps
      -- 
    sendModule_CP_7961_elements(72) <= sendModule_CP_7961_elements(73);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	72 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3212_update_completed_
      -- 
    -- Element group sendModule_CP_7961_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => sendModule_CP_7961_elements(71), ack => sendModule_CP_7961_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_sample_start__ps
      -- CP-element group 74: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_Sample/req
      -- 
    req_8174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(74), ack => n_chl_3268_3213_buf_req_0); -- 
    -- Element group sendModule_CP_7961_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_update_start__ps
      -- CP-element group 75: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_update_start_
      -- CP-element group 75: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_Update/req
      -- 
    req_8179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(75), ack => n_chl_3268_3213_buf_req_1); -- 
    -- Element group sendModule_CP_7961_elements(75) is bound as output of CP function.
    -- CP-element group 76:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_Sample/ack
      -- 
    ack_8175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3268_3213_buf_ack_0, ack => sendModule_CP_7961_elements(76)); -- 
    -- CP-element group 77:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_Update/ack
      -- CP-element group 77: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_chl_3213_Update/$exit
      -- 
    ack_8180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3268_3213_buf_ack_1, ack => sendModule_CP_7961_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	15 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	18 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	17 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_sample_start_
      -- 
    sendModule_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(18);
      gj_sendModule_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	15 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	19 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_update_start_
      -- 
    sendModule_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(83);
      gj_sendModule_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_sample_start__ps
      -- 
    sendModule_CP_7961_elements(80) <= sendModule_CP_7961_elements(17);
    -- CP-element group 81:  join  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	18 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7961_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	19 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_update_start__ps
      -- 
    sendModule_CP_7961_elements(82) <= sendModule_CP_7961_elements(19);
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	20 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_update_completed__ps
      -- 
    -- Element group sendModule_CP_7961_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	13 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_loopback_trigger
      -- 
    sendModule_CP_7961_elements(84) <= sendModule_CP_7961_elements(13);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_loopback_sample_req_ps
      -- CP-element group 85: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_loopback_sample_req
      -- 
    phi_stmt_3214_loopback_sample_req_8191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3214_loopback_sample_req_8191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(85), ack => phi_stmt_3214_req_1); -- 
    -- Element group sendModule_CP_7961_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	14 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_entry_trigger
      -- 
    sendModule_CP_7961_elements(86) <= sendModule_CP_7961_elements(14);
    -- CP-element group 87:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_entry_sample_req
      -- CP-element group 87: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_entry_sample_req_ps
      -- 
    phi_stmt_3214_entry_sample_req_8194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3214_entry_sample_req_8194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(87), ack => phi_stmt_3214_req_0); -- 
    -- Element group sendModule_CP_7961_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_phi_mux_ack
      -- CP-element group 88: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3214_phi_mux_ack_ps
      -- 
    phi_stmt_3214_phi_mux_ack_8197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3214_ack_0, ack => sendModule_CP_7961_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3217_sample_start__ps
      -- CP-element group 89: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3217_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3217_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3217_sample_completed_
      -- 
    -- Element group sendModule_CP_7961_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3217_update_start__ps
      -- CP-element group 90: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3217_update_start_
      -- 
    -- Element group sendModule_CP_7961_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3217_update_completed__ps
      -- 
    sendModule_CP_7961_elements(91) <= sendModule_CP_7961_elements(92);
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3217_update_completed_
      -- 
    -- Element group sendModule_CP_7961_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => sendModule_CP_7961_elements(90), ack => sendModule_CP_7961_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_Sample/req
      -- CP-element group 93: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_sample_start__ps
      -- 
    req_8218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(93), ack => n_col_3249_3218_buf_req_0); -- 
    -- Element group sendModule_CP_7961_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_update_start_
      -- CP-element group 94: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_update_start__ps
      -- CP-element group 94: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_Update/req
      -- CP-element group 94: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_Update/$entry
      -- 
    req_8223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(94), ack => n_col_3249_3218_buf_req_1); -- 
    -- Element group sendModule_CP_7961_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_Sample/ack
      -- CP-element group 95: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_sample_completed__ps
      -- 
    ack_8219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3249_3218_buf_ack_0, ack => sendModule_CP_7961_elements(95)); -- 
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_Update/ack
      -- CP-element group 96: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_col_3218_Update/$exit
      -- 
    ack_8224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3249_3218_buf_ack_1, ack => sendModule_CP_7961_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	15 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	119 
    -- CP-element group 97: 	18 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	17 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_sample_start_
      -- 
    sendModule_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(119) & sendModule_CP_7961_elements(18);
      gj_sendModule_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	15 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	19 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_update_start_
      -- 
    sendModule_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(102);
      gj_sendModule_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	17 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_sample_start__ps
      -- 
    sendModule_CP_7961_elements(99) <= sendModule_CP_7961_elements(17);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	18 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_sample_completed__ps
      -- 
    -- Element group sendModule_CP_7961_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	19 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_update_start__ps
      -- 
    sendModule_CP_7961_elements(101) <= sendModule_CP_7961_elements(19);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	20 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_update_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_update_completed_
      -- 
    -- Element group sendModule_CP_7961_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	13 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_loopback_trigger
      -- 
    sendModule_CP_7961_elements(103) <= sendModule_CP_7961_elements(13);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_loopback_sample_req_ps
      -- CP-element group 104: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_loopback_sample_req
      -- 
    phi_stmt_3219_loopback_sample_req_8235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3219_loopback_sample_req_8235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(104), ack => phi_stmt_3219_req_1); -- 
    -- Element group sendModule_CP_7961_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	14 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_entry_trigger
      -- 
    sendModule_CP_7961_elements(105) <= sendModule_CP_7961_elements(14);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_entry_sample_req_ps
      -- CP-element group 106: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_entry_sample_req
      -- 
    phi_stmt_3219_entry_sample_req_8238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3219_entry_sample_req_8238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(106), ack => phi_stmt_3219_req_0); -- 
    -- Element group sendModule_CP_7961_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_phi_mux_ack_ps
      -- CP-element group 107: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/phi_stmt_3219_phi_mux_ack
      -- 
    phi_stmt_3219_phi_mux_ack_8241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3219_ack_0, ack => sendModule_CP_7961_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3222_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3222_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3222_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3222_sample_start__ps
      -- 
    -- Element group sendModule_CP_7961_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3222_update_start_
      -- CP-element group 109: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3222_update_start__ps
      -- 
    -- Element group sendModule_CP_7961_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3222_update_completed__ps
      -- 
    sendModule_CP_7961_elements(110) <= sendModule_CP_7961_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3222_update_completed_
      -- 
    -- Element group sendModule_CP_7961_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => sendModule_CP_7961_elements(109), ack => sendModule_CP_7961_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_Sample/req
      -- CP-element group 112: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_sample_start__ps
      -- 
    req_8262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(112), ack => n_row_3260_3223_buf_req_0); -- 
    -- Element group sendModule_CP_7961_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_Update/req
      -- CP-element group 113: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_update_start_
      -- CP-element group 113: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_update_start__ps
      -- 
    req_8267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(113), ack => n_row_3260_3223_buf_req_1); -- 
    -- Element group sendModule_CP_7961_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_sample_completed__ps
      -- 
    ack_8263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3260_3223_buf_ack_0, ack => sendModule_CP_7961_elements(114)); -- 
    -- CP-element group 115:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_Update/ack
      -- CP-element group 115: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/R_n_row_3223_update_completed__ps
      -- 
    ack_8268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3260_3223_buf_ack_1, ack => sendModule_CP_7961_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	15 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_sample_start_
      -- 
    rr_8277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(116), ack => SUB_u16_u16_3233_inst_req_0); -- 
    sendModule_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(118);
      gj_sendModule_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	18 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_update_start_
      -- CP-element group 117: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_Update/cr
      -- 
    cr_8282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(117), ack => SUB_u16_u16_3233_inst_req_1); -- 
    sendModule_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(18) & sendModule_CP_7961_elements(119);
      gj_sendModule_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_sample_completed_
      -- 
    ra_8278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3233_inst_ack_0, ack => sendModule_CP_7961_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	16 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	21 
    -- CP-element group 119: 	38 
    -- CP-element group 119: 	59 
    -- CP-element group 119: 	97 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3233_Update/$exit
      -- 
    ca_8283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3233_inst_ack_1, ack => sendModule_CP_7961_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	15 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_sample_start_
      -- 
    rr_8291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(120), ack => type_cast_3271_inst_req_0); -- 
    sendModule_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(122);
      gj_sendModule_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	18 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_update_start_
      -- 
    cr_8296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(121), ack => type_cast_3271_inst_req_1); -- 
    sendModule_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(18) & sendModule_CP_7961_elements(123);
      gj_sendModule_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_sample_completed_
      -- 
    ra_8292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3271_inst_ack_0, ack => sendModule_CP_7961_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	286 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	21 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3271_update_completed_
      -- 
    ca_8297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3271_inst_ack_1, ack => sendModule_CP_7961_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	15 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_Sample/rr
      -- 
    rr_8305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(124), ack => type_cast_3280_inst_req_0); -- 
    sendModule_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(126);
      gj_sendModule_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	18 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_update_start_
      -- CP-element group 125: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_Update/cr
      -- CP-element group 125: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_Update/$entry
      -- 
    cr_8310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(125), ack => type_cast_3280_inst_req_1); -- 
    sendModule_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(18) & sendModule_CP_7961_elements(127);
      gj_sendModule_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_Sample/ra
      -- 
    ra_8306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3280_inst_ack_0, ack => sendModule_CP_7961_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	286 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	38 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/type_cast_3280_Update/$exit
      -- 
    ca_8311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3280_inst_ack_1, ack => sendModule_CP_7961_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	132 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	133 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_request/$entry
      -- CP-element group 128: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_request/req
      -- 
    req_8351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(128), ack => addr_of_3321_final_reg_req_0); -- 
    sendModule_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(132) & sendModule_CP_7961_elements(133);
      gj_sendModule_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	15 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	256 
    -- CP-element group 129: 	144 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	134 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_update_start_
      -- CP-element group 129: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_complete/req
      -- CP-element group 129: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_complete/$entry
      -- 
    req_8356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(129), ack => addr_of_3321_final_reg_req_1); -- 
    sendModule_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(256) & sendModule_CP_7961_elements(144);
      gj_sendModule_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	15 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	133 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_update_start
      -- CP-element group 130: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_Update/req
      -- CP-element group 130: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_Update/$entry
      -- 
    req_8341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(130), ack => array_obj_ref_3320_index_offset_req_1); -- 
    sendModule_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(133);
      gj_sendModule_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	24 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	286 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	22 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_sample_complete
      -- CP-element group 131: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_Sample/ack
      -- CP-element group 131: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_Sample/$exit
      -- 
    ack_8337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3320_index_offset_ack_0, ack => sendModule_CP_7961_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	128 
    -- CP-element group 132:  members (8) 
      -- CP-element group 132: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_base_plus_offset/sum_rename_req
      -- CP-element group 132: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_root_address_calculated
      -- CP-element group 132: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_offset_calculated
      -- CP-element group 132: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_base_plus_offset/sum_rename_ack
      -- CP-element group 132: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_base_plus_offset/$exit
      -- CP-element group 132: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_base_plus_offset/$entry
      -- CP-element group 132: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_Update/ack
      -- CP-element group 132: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3320_final_index_sum_regn_Update/$exit
      -- 
    ack_8342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3320_index_offset_ack_1, ack => sendModule_CP_7961_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: 	128 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_request/ack
      -- CP-element group 133: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_request/$exit
      -- 
    ack_8352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3321_final_reg_ack_0, ack => sendModule_CP_7961_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	129 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	142 
    -- CP-element group 134: 	254 
    -- CP-element group 134:  members (19) 
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_plus_offset/sum_rename_req
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_word_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_plus_offset/sum_rename_ack
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_addr_resize/base_resize_req
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_root_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_addr_resize/$exit
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_word_addrgen/$entry
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_address_resized
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_plus_offset/$exit
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_plus_offset/$entry
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_addr_resize/base_resize_ack
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_word_addrgen/root_register_ack
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_word_addrgen/root_register_req
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_word_addrgen/$exit
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_base_addr_resize/$entry
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_complete/ack
      -- CP-element group 134: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3321_complete/$exit
      -- 
    ack_8357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3321_final_reg_ack_1, ack => sendModule_CP_7961_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	139 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	140 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	140 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_request/req
      -- CP-element group 135: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_request/$entry
      -- 
    req_8397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(135), ack => addr_of_3331_final_reg_req_0); -- 
    sendModule_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(139) & sendModule_CP_7961_elements(140);
      gj_sendModule_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	15 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	148 
    -- CP-element group 136: 	268 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	141 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_complete/req
      -- CP-element group 136: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_update_start_
      -- 
    req_8402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(136), ack => addr_of_3331_final_reg_req_1); -- 
    sendModule_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(148) & sendModule_CP_7961_elements(268);
      gj_sendModule_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	15 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	140 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_Update/req
      -- CP-element group 137: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_update_start
      -- 
    req_8387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(137), ack => array_obj_ref_3330_index_offset_req_1); -- 
    sendModule_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(140);
      gj_sendModule_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	43 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	286 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	39 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_sample_complete
      -- CP-element group 138: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_Sample/ack
      -- 
    ack_8383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3330_index_offset_ack_0, ack => sendModule_CP_7961_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	135 
    -- CP-element group 139:  members (8) 
      -- CP-element group 139: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_base_plus_offset/$exit
      -- CP-element group 139: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_base_plus_offset/sum_rename_req
      -- CP-element group 139: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_final_index_sum_regn_Update/ack
      -- CP-element group 139: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_base_plus_offset/$entry
      -- CP-element group 139: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_base_plus_offset/sum_rename_ack
      -- CP-element group 139: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_offset_calculated
      -- CP-element group 139: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/array_obj_ref_3330_root_address_calculated
      -- 
    ack_8388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3330_index_offset_ack_1, ack => sendModule_CP_7961_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	135 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	135 
    -- CP-element group 140: 	137 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_request/ack
      -- CP-element group 140: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_request/$exit
      -- 
    ack_8398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3331_final_reg_ack_0, ack => sendModule_CP_7961_elements(140)); -- 
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	136 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	266 
    -- CP-element group 141: 	146 
    -- CP-element group 141:  members (19) 
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_addr_resize/base_resize_req
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_address_resized
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_word_addrgen/$exit
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_word_addrgen/$entry
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_addr_resize/base_resize_ack
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_word_addrgen/root_register_ack
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_addr_resize/$entry
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_addr_resize/$exit
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_word_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_word_addrgen/root_register_req
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_complete/ack
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_complete/$exit
      -- CP-element group 141: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/addr_of_3331_update_completed_
      -- 
    ack_8403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3331_final_reg_ack_1, ack => sendModule_CP_7961_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	134 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	276 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (5) 
      -- CP-element group 142: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Sample/word_access_start/word_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Sample/word_access_start/word_0/rr
      -- CP-element group 142: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Sample/word_access_start/$entry
      -- CP-element group 142: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_sample_start_
      -- 
    rr_8436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(142), ack => ptr_deref_3335_load_0_req_0); -- 
    sendModule_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(134) & sendModule_CP_7961_elements(276);
      gj_sendModule_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	168 
    -- CP-element group 143: 	172 
    -- CP-element group 143: 	160 
    -- CP-element group 143: 	164 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/word_access_complete/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/word_access_complete/$entry
      -- CP-element group 143: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/word_access_complete/word_0/cr
      -- CP-element group 143: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_update_start_
      -- 
    cr_8447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(143), ack => ptr_deref_3335_load_0_req_1); -- 
    sendModule_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(168) & sendModule_CP_7961_elements(172) & sendModule_CP_7961_elements(160) & sendModule_CP_7961_elements(164);
      gj_sendModule_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	283 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	129 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Sample/word_access_start/word_0/ra
      -- CP-element group 144: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_sample_completed_
      -- 
    ra_8437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3335_load_0_ack_0, ack => sendModule_CP_7961_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	170 
    -- CP-element group 145: 	158 
    -- CP-element group 145: 	162 
    -- CP-element group 145: 	166 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/ptr_deref_3335_Merge/$entry
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/ptr_deref_3335_Merge/$exit
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/ptr_deref_3335_Merge/merge_ack
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/ptr_deref_3335_Merge/merge_req
      -- CP-element group 145: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_Update/word_access_complete/word_0/ca
      -- 
    ca_8448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3335_load_0_ack_1, ack => sendModule_CP_7961_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	141 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	276 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Sample/word_access_start/$entry
      -- CP-element group 146: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Sample/word_access_start/word_0/rr
      -- CP-element group 146: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Sample/word_access_start/word_0/$entry
      -- 
    rr_8486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(146), ack => ptr_deref_3339_load_0_req_0); -- 
    sendModule_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(141) & sendModule_CP_7961_elements(276);
      gj_sendModule_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	180 
    -- CP-element group 147: 	184 
    -- CP-element group 147: 	188 
    -- CP-element group 147: 	176 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/word_access_complete/word_0/cr
      -- CP-element group 147: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_update_start_
      -- CP-element group 147: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/word_access_complete/word_0/$entry
      -- CP-element group 147: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/word_access_complete/$entry
      -- 
    cr_8497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(147), ack => ptr_deref_3339_load_0_req_1); -- 
    sendModule_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(180) & sendModule_CP_7961_elements(184) & sendModule_CP_7961_elements(188) & sendModule_CP_7961_elements(176);
      gj_sendModule_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	284 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	136 
    -- CP-element group 148:  members (5) 
      -- CP-element group 148: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Sample/word_access_start/$exit
      -- CP-element group 148: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Sample/word_access_start/word_0/ra
      -- CP-element group 148: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Sample/word_access_start/word_0/$exit
      -- 
    ra_8487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3339_load_0_ack_0, ack => sendModule_CP_7961_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	182 
    -- CP-element group 149: 	186 
    -- CP-element group 149: 	174 
    -- CP-element group 149: 	178 
    -- CP-element group 149:  members (9) 
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/word_access_complete/word_0/ca
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/ptr_deref_3339_Merge/$entry
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/ptr_deref_3339_Merge/$exit
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/word_access_complete/word_0/$exit
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/ptr_deref_3339_Merge/merge_req
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/ptr_deref_3339_Merge/merge_ack
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_Update/word_access_complete/$exit
      -- CP-element group 149: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_update_completed_
      -- 
    ca_8498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3339_load_0_ack_1, ack => sendModule_CP_7961_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	15 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_Sample/$entry
      -- 
    rr_8511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(150), ack => RPIPE_output_pipe_3342_inst_req_0); -- 
    sendModule_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(153);
      gj_sendModule_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	212 
    -- CP-element group 151: 	220 
    -- CP-element group 151: 	196 
    -- CP-element group 151: 	204 
    -- CP-element group 151: 	157 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_Update/cr
      -- CP-element group 151: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_update_start_
      -- 
    cr_8516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(151), ack => RPIPE_output_pipe_3342_inst_req_1); -- 
    sendModule_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(152) & sendModule_CP_7961_elements(212) & sendModule_CP_7961_elements(220) & sendModule_CP_7961_elements(196) & sendModule_CP_7961_elements(204) & sendModule_CP_7961_elements(157);
      gj_sendModule_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	151 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_Sample/$exit
      -- 
    ra_8512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3342_inst_ack_0, ack => sendModule_CP_7961_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	210 
    -- CP-element group 153: 	218 
    -- CP-element group 153: 	194 
    -- CP-element group 153: 	202 
    -- CP-element group 153: 	154 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3342_update_completed_
      -- 
    ca_8517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3342_inst_ack_1, ack => sendModule_CP_7961_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	157 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_Sample/rr
      -- 
    rr_8525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(154), ack => RPIPE_output_pipe_3345_inst_req_0); -- 
    sendModule_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(153) & sendModule_CP_7961_elements(157);
      gj_sendModule_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	252 
    -- CP-element group 155: 	236 
    -- CP-element group 155: 	244 
    -- CP-element group 155: 	228 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_update_start_
      -- CP-element group 155: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_Update/cr
      -- 
    cr_8530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(155), ack => RPIPE_output_pipe_3345_inst_req_1); -- 
    sendModule_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(156) & sendModule_CP_7961_elements(252) & sendModule_CP_7961_elements(236) & sendModule_CP_7961_elements(244) & sendModule_CP_7961_elements(228);
      gj_sendModule_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	155 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_Sample/ra
      -- 
    ra_8526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3345_inst_ack_0, ack => sendModule_CP_7961_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	250 
    -- CP-element group 157: 	242 
    -- CP-element group 157: 	226 
    -- CP-element group 157: 	234 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	151 
    -- CP-element group 157: 	154 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/RPIPE_output_pipe_3345_Update/ca
      -- 
    ca_8531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3345_inst_ack_1, ack => sendModule_CP_7961_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	145 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_Sample/rr
      -- 
    rr_8539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(158), ack => slice_3349_inst_req_0); -- 
    sendModule_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(145) & sendModule_CP_7961_elements(160);
      gj_sendModule_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	260 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_update_start_
      -- CP-element group 159: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_Update/cr
      -- 
    cr_8544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(159), ack => slice_3349_inst_req_1); -- 
    sendModule_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	143 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_Sample/ra
      -- 
    ra_8540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3349_inst_ack_0, ack => sendModule_CP_7961_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	258 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3349_Update/ca
      -- 
    ca_8545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3349_inst_ack_1, ack => sendModule_CP_7961_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	145 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_Sample/rr
      -- 
    rr_8553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(162), ack => slice_3353_inst_req_0); -- 
    sendModule_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(145) & sendModule_CP_7961_elements(164);
      gj_sendModule_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	260 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_Update/cr
      -- 
    cr_8558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(163), ack => slice_3353_inst_req_1); -- 
    sendModule_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	143 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_Sample/ra
      -- 
    ra_8554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3353_inst_ack_0, ack => sendModule_CP_7961_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	258 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3353_Update/ca
      -- 
    ca_8559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3353_inst_ack_1, ack => sendModule_CP_7961_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	145 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_Sample/rr
      -- 
    rr_8567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(166), ack => slice_3357_inst_req_0); -- 
    sendModule_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(145) & sendModule_CP_7961_elements(168);
      gj_sendModule_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	260 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_update_start_
      -- CP-element group 167: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_Update/cr
      -- 
    cr_8572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(167), ack => slice_3357_inst_req_1); -- 
    sendModule_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	143 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_Sample/ra
      -- 
    ra_8568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3357_inst_ack_0, ack => sendModule_CP_7961_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	258 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3357_Update/ca
      -- 
    ca_8573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3357_inst_ack_1, ack => sendModule_CP_7961_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	145 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_Sample/rr
      -- 
    rr_8581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(170), ack => slice_3361_inst_req_0); -- 
    sendModule_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(145) & sendModule_CP_7961_elements(172);
      gj_sendModule_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	260 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_update_start_
      -- CP-element group 171: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_Update/cr
      -- 
    cr_8586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(171), ack => slice_3361_inst_req_1); -- 
    sendModule_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	143 
    -- CP-element group 172: 	170 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_Sample/ra
      -- 
    ra_8582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3361_inst_ack_0, ack => sendModule_CP_7961_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	258 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3361_Update/ca
      -- 
    ca_8587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3361_inst_ack_1, ack => sendModule_CP_7961_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	149 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_Sample/rr
      -- 
    rr_8595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(174), ack => slice_3365_inst_req_0); -- 
    sendModule_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(149) & sendModule_CP_7961_elements(176);
      gj_sendModule_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	272 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_update_start_
      -- CP-element group 175: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_Update/cr
      -- 
    cr_8600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(175), ack => slice_3365_inst_req_1); -- 
    sendModule_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: 	147 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_Sample/ra
      -- 
    ra_8596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3365_inst_ack_0, ack => sendModule_CP_7961_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	270 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3365_Update/ca
      -- 
    ca_8601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3365_inst_ack_1, ack => sendModule_CP_7961_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	149 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_Sample/rr
      -- 
    rr_8609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(178), ack => slice_3369_inst_req_0); -- 
    sendModule_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(149) & sendModule_CP_7961_elements(180);
      gj_sendModule_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	272 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_update_start_
      -- CP-element group 179: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_Update/cr
      -- 
    cr_8614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(179), ack => slice_3369_inst_req_1); -- 
    sendModule_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: 	147 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_Sample/ra
      -- 
    ra_8610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3369_inst_ack_0, ack => sendModule_CP_7961_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	270 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3369_Update/ca
      -- 
    ca_8615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3369_inst_ack_1, ack => sendModule_CP_7961_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	149 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_Sample/rr
      -- 
    rr_8623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(182), ack => slice_3373_inst_req_0); -- 
    sendModule_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(149) & sendModule_CP_7961_elements(184);
      gj_sendModule_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	272 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_update_start_
      -- CP-element group 183: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_Update/cr
      -- 
    cr_8628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(183), ack => slice_3373_inst_req_1); -- 
    sendModule_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	147 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_Sample/ra
      -- 
    ra_8624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3373_inst_ack_0, ack => sendModule_CP_7961_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	270 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3373_Update/ca
      -- 
    ca_8629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3373_inst_ack_1, ack => sendModule_CP_7961_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	149 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_Sample/rr
      -- 
    rr_8637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(186), ack => slice_3377_inst_req_0); -- 
    sendModule_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(149) & sendModule_CP_7961_elements(188);
      gj_sendModule_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	272 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_update_start_
      -- CP-element group 187: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_Update/cr
      -- 
    cr_8642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(187), ack => slice_3377_inst_req_1); -- 
    sendModule_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: 	147 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_Sample/ra
      -- 
    ra_8638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3377_inst_ack_0, ack => sendModule_CP_7961_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	270 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/slice_3377_Update/ca
      -- 
    ca_8643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3377_inst_ack_1, ack => sendModule_CP_7961_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	24 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_Sample/rr
      -- 
    rr_8651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(190), ack => EQ_u2_u1_3390_inst_req_0); -- 
    sendModule_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(24) & sendModule_CP_7961_elements(192);
      gj_sendModule_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	260 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_update_start_
      -- CP-element group 191: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_Update/cr
      -- 
    cr_8656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(191), ack => EQ_u2_u1_3390_inst_req_1); -- 
    sendModule_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	22 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_Sample/ra
      -- 
    ra_8652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3390_inst_ack_0, ack => sendModule_CP_7961_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	258 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3390_Update/ca
      -- 
    ca_8657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3390_inst_ack_1, ack => sendModule_CP_7961_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	153 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_Sample/req
      -- 
    req_8665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(194), ack => W_output_data1_3262_delayed_14_0_3392_inst_req_0); -- 
    sendModule_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(153) & sendModule_CP_7961_elements(196);
      gj_sendModule_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	260 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_update_start_
      -- CP-element group 195: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_Update/req
      -- 
    req_8670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(195), ack => W_output_data1_3262_delayed_14_0_3392_inst_req_1); -- 
    sendModule_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	151 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_Sample/ack
      -- 
    ack_8666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3262_delayed_14_0_3392_inst_ack_0, ack => sendModule_CP_7961_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	258 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3394_Update/ack
      -- 
    ack_8671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3262_delayed_14_0_3392_inst_ack_1, ack => sendModule_CP_7961_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	24 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_Sample/rr
      -- 
    rr_8679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(198), ack => EQ_u2_u1_3404_inst_req_0); -- 
    sendModule_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(24) & sendModule_CP_7961_elements(200);
      gj_sendModule_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	260 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_update_start_
      -- CP-element group 199: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_Update/cr
      -- 
    cr_8684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(199), ack => EQ_u2_u1_3404_inst_req_1); -- 
    sendModule_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	22 
    -- CP-element group 200: 	198 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_Sample/ra
      -- 
    ra_8680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3404_inst_ack_0, ack => sendModule_CP_7961_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	258 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3404_Update/ca
      -- 
    ca_8685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3404_inst_ack_1, ack => sendModule_CP_7961_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	153 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_Sample/req
      -- 
    req_8693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(202), ack => W_output_data1_3270_delayed_14_0_3406_inst_req_0); -- 
    sendModule_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(153) & sendModule_CP_7961_elements(204);
      gj_sendModule_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	260 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_update_start_
      -- CP-element group 203: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_Update/req
      -- 
    req_8698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(203), ack => W_output_data1_3270_delayed_14_0_3406_inst_req_1); -- 
    sendModule_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	151 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_Sample/ack
      -- 
    ack_8694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3270_delayed_14_0_3406_inst_ack_0, ack => sendModule_CP_7961_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	258 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3408_Update/ack
      -- 
    ack_8699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3270_delayed_14_0_3406_inst_ack_1, ack => sendModule_CP_7961_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	24 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_Sample/rr
      -- 
    rr_8707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(206), ack => EQ_u2_u1_3418_inst_req_0); -- 
    sendModule_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(24) & sendModule_CP_7961_elements(208);
      gj_sendModule_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	260 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_update_start_
      -- CP-element group 207: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_Update/cr
      -- 
    cr_8712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(207), ack => EQ_u2_u1_3418_inst_req_1); -- 
    sendModule_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	22 
    -- CP-element group 208: 	206 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_Sample/ra
      -- 
    ra_8708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3418_inst_ack_0, ack => sendModule_CP_7961_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	258 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3418_Update/ca
      -- 
    ca_8713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3418_inst_ack_1, ack => sendModule_CP_7961_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	153 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_Sample/req
      -- 
    req_8721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(210), ack => W_output_data1_3278_delayed_14_0_3420_inst_req_0); -- 
    sendModule_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(153) & sendModule_CP_7961_elements(212);
      gj_sendModule_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	260 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_update_start_
      -- CP-element group 211: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_Update/req
      -- 
    req_8726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(211), ack => W_output_data1_3278_delayed_14_0_3420_inst_req_1); -- 
    sendModule_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	151 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_Sample/ack
      -- 
    ack_8722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3278_delayed_14_0_3420_inst_ack_0, ack => sendModule_CP_7961_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	258 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3422_Update/ack
      -- 
    ack_8727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3278_delayed_14_0_3420_inst_ack_1, ack => sendModule_CP_7961_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	24 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_Sample/rr
      -- 
    rr_8735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(214), ack => EQ_u2_u1_3432_inst_req_0); -- 
    sendModule_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(24) & sendModule_CP_7961_elements(216);
      gj_sendModule_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	260 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_update_start_
      -- CP-element group 215: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_Update/cr
      -- 
    cr_8740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(215), ack => EQ_u2_u1_3432_inst_req_1); -- 
    sendModule_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	22 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_Sample/ra
      -- 
    ra_8736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3432_inst_ack_0, ack => sendModule_CP_7961_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	258 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3432_Update/ca
      -- 
    ca_8741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3432_inst_ack_1, ack => sendModule_CP_7961_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	153 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_Sample/req
      -- 
    req_8749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(218), ack => W_output_data1_3286_delayed_14_0_3434_inst_req_0); -- 
    sendModule_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(153) & sendModule_CP_7961_elements(220);
      gj_sendModule_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	260 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_update_start_
      -- CP-element group 219: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_Update/req
      -- 
    req_8754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(219), ack => W_output_data1_3286_delayed_14_0_3434_inst_req_1); -- 
    sendModule_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	151 
    -- CP-element group 220: 	218 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_Sample/ack
      -- 
    ack_8750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3286_delayed_14_0_3434_inst_ack_0, ack => sendModule_CP_7961_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	258 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3436_Update/ack
      -- 
    ack_8755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3286_delayed_14_0_3434_inst_ack_1, ack => sendModule_CP_7961_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	43 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_Sample/rr
      -- 
    rr_8763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(222), ack => EQ_u2_u1_3446_inst_req_0); -- 
    sendModule_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(43) & sendModule_CP_7961_elements(224);
      gj_sendModule_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	272 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_update_start_
      -- CP-element group 223: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_Update/cr
      -- 
    cr_8768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(223), ack => EQ_u2_u1_3446_inst_req_1); -- 
    sendModule_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: 	39 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_Sample/ra
      -- 
    ra_8764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3446_inst_ack_0, ack => sendModule_CP_7961_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	270 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3446_Update/ca
      -- 
    ca_8769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3446_inst_ack_1, ack => sendModule_CP_7961_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	157 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_Sample/req
      -- 
    req_8777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(226), ack => W_output_data2_3294_delayed_14_0_3448_inst_req_0); -- 
    sendModule_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(157) & sendModule_CP_7961_elements(228);
      gj_sendModule_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	272 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_update_start_
      -- CP-element group 227: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_Update/req
      -- 
    req_8782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(227), ack => W_output_data2_3294_delayed_14_0_3448_inst_req_1); -- 
    sendModule_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: 	155 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_Sample/ack
      -- 
    ack_8778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3294_delayed_14_0_3448_inst_ack_0, ack => sendModule_CP_7961_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	270 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3450_Update/ack
      -- 
    ack_8783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3294_delayed_14_0_3448_inst_ack_1, ack => sendModule_CP_7961_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	43 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_Sample/rr
      -- 
    rr_8791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(230), ack => EQ_u2_u1_3460_inst_req_0); -- 
    sendModule_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(43) & sendModule_CP_7961_elements(232);
      gj_sendModule_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	272 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	233 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_update_start_
      -- CP-element group 231: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_Update/cr
      -- 
    cr_8796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(231), ack => EQ_u2_u1_3460_inst_req_1); -- 
    sendModule_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: 	39 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_Sample/ra
      -- 
    ra_8792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3460_inst_ack_0, ack => sendModule_CP_7961_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	270 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3460_Update/ca
      -- 
    ca_8797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3460_inst_ack_1, ack => sendModule_CP_7961_elements(233)); -- 
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	157 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_Sample/req
      -- 
    req_8805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(234), ack => W_output_data2_3302_delayed_14_0_3462_inst_req_0); -- 
    sendModule_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(157) & sendModule_CP_7961_elements(236);
      gj_sendModule_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: marked-predecessors 
    -- CP-element group 235: 	272 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_update_start_
      -- CP-element group 235: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_Update/req
      -- 
    req_8810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(235), ack => W_output_data2_3302_delayed_14_0_3462_inst_req_1); -- 
    sendModule_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	155 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_Sample/ack
      -- 
    ack_8806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3302_delayed_14_0_3462_inst_ack_0, ack => sendModule_CP_7961_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	270 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3464_Update/ack
      -- 
    ack_8811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3302_delayed_14_0_3462_inst_ack_1, ack => sendModule_CP_7961_elements(237)); -- 
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	43 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_Sample/rr
      -- 
    rr_8819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(238), ack => EQ_u2_u1_3474_inst_req_0); -- 
    sendModule_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(43) & sendModule_CP_7961_elements(240);
      gj_sendModule_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: marked-predecessors 
    -- CP-element group 239: 	272 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_update_start_
      -- CP-element group 239: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_Update/cr
      -- 
    cr_8824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(239), ack => EQ_u2_u1_3474_inst_req_1); -- 
    sendModule_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: 	39 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_Sample/ra
      -- 
    ra_8820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3474_inst_ack_0, ack => sendModule_CP_7961_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	270 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3474_Update/ca
      -- 
    ca_8825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3474_inst_ack_1, ack => sendModule_CP_7961_elements(241)); -- 
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	157 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_Sample/req
      -- 
    req_8833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(242), ack => W_output_data2_3310_delayed_14_0_3476_inst_req_0); -- 
    sendModule_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(157) & sendModule_CP_7961_elements(244);
      gj_sendModule_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: marked-predecessors 
    -- CP-element group 243: 	272 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	245 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_update_start_
      -- CP-element group 243: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_Update/req
      -- 
    req_8838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(243), ack => W_output_data2_3310_delayed_14_0_3476_inst_req_1); -- 
    sendModule_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	155 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_Sample/ack
      -- 
    ack_8834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3310_delayed_14_0_3476_inst_ack_0, ack => sendModule_CP_7961_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	243 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	270 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3478_Update/ack
      -- 
    ack_8839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3310_delayed_14_0_3476_inst_ack_1, ack => sendModule_CP_7961_elements(245)); -- 
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	43 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_Sample/rr
      -- 
    rr_8847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(246), ack => EQ_u2_u1_3488_inst_req_0); -- 
    sendModule_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(43) & sendModule_CP_7961_elements(248);
      gj_sendModule_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: marked-predecessors 
    -- CP-element group 247: 	272 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_update_start_
      -- CP-element group 247: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_Update/cr
      -- 
    cr_8852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(247), ack => EQ_u2_u1_3488_inst_req_1); -- 
    sendModule_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: 	39 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_Sample/ra
      -- 
    ra_8848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3488_inst_ack_0, ack => sendModule_CP_7961_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	270 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/EQ_u2_u1_3488_Update/ca
      -- 
    ca_8853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u2_u1_3488_inst_ack_1, ack => sendModule_CP_7961_elements(249)); -- 
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	157 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_Sample/req
      -- 
    req_8861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(250), ack => W_output_data2_3318_delayed_14_0_3490_inst_req_0); -- 
    sendModule_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(157) & sendModule_CP_7961_elements(252);
      gj_sendModule_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: marked-predecessors 
    -- CP-element group 251: 	272 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_update_start_
      -- CP-element group 251: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_Update/req
      -- 
    req_8866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(251), ack => W_output_data2_3318_delayed_14_0_3490_inst_req_1); -- 
    sendModule_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	155 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_Sample/ack
      -- 
    ack_8862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3318_delayed_14_0_3490_inst_ack_0, ack => sendModule_CP_7961_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	270 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3492_Update/ack
      -- 
    ack_8867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3318_delayed_14_0_3490_inst_ack_1, ack => sendModule_CP_7961_elements(253)); -- 
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	134 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_Sample/req
      -- 
    req_8875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(254), ack => W_fetch_addr1_3322_delayed_8_0_3499_inst_req_0); -- 
    sendModule_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(134) & sendModule_CP_7961_elements(256);
      gj_sendModule_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: marked-predecessors 
    -- CP-element group 255: 	264 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_update_start_
      -- CP-element group 255: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_Update/req
      -- 
    req_8880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(255), ack => W_fetch_addr1_3322_delayed_8_0_3499_inst_req_1); -- 
    sendModule_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(264);
      gj_sendModule_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	129 
    -- CP-element group 256: 	254 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_Sample/ack
      -- 
    ack_8876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr1_3322_delayed_8_0_3499_inst_ack_0, ack => sendModule_CP_7961_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	262 
    -- CP-element group 257:  members (19) 
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3501_Update/ack
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_address_calculated
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_word_address_calculated
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_root_address_calculated
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_address_resized
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_addr_resize/$entry
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_addr_resize/$exit
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_addr_resize/base_resize_req
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_addr_resize/base_resize_ack
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_plus_offset/$entry
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_plus_offset/$exit
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_plus_offset/sum_rename_req
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_base_plus_offset/sum_rename_ack
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_word_addrgen/$entry
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_word_addrgen/$exit
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_word_addrgen/root_register_req
      -- CP-element group 257: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_word_addrgen/root_register_ack
      -- 
    ack_8881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr1_3322_delayed_8_0_3499_inst_ack_1, ack => sendModule_CP_7961_elements(257)); -- 
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	209 
    -- CP-element group 258: 	213 
    -- CP-element group 258: 	217 
    -- CP-element group 258: 	221 
    -- CP-element group 258: 	197 
    -- CP-element group 258: 	201 
    -- CP-element group 258: 	205 
    -- CP-element group 258: 	193 
    -- CP-element group 258: 	169 
    -- CP-element group 258: 	173 
    -- CP-element group 258: 	161 
    -- CP-element group 258: 	165 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_Sample/rr
      -- 
    rr_8889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(258), ack => CONCAT_u32_u64_3510_inst_req_0); -- 
    sendModule_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(209) & sendModule_CP_7961_elements(213) & sendModule_CP_7961_elements(217) & sendModule_CP_7961_elements(221) & sendModule_CP_7961_elements(197) & sendModule_CP_7961_elements(201) & sendModule_CP_7961_elements(205) & sendModule_CP_7961_elements(193) & sendModule_CP_7961_elements(169) & sendModule_CP_7961_elements(173) & sendModule_CP_7961_elements(161) & sendModule_CP_7961_elements(165) & sendModule_CP_7961_elements(260);
      gj_sendModule_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: marked-predecessors 
    -- CP-element group 259: 	264 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	261 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_update_start_
      -- CP-element group 259: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_Update/cr
      -- 
    cr_8894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(259), ack => CONCAT_u32_u64_3510_inst_req_1); -- 
    sendModule_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(264);
      gj_sendModule_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	211 
    -- CP-element group 260: 	215 
    -- CP-element group 260: 	219 
    -- CP-element group 260: 	195 
    -- CP-element group 260: 	199 
    -- CP-element group 260: 	203 
    -- CP-element group 260: 	207 
    -- CP-element group 260: 	191 
    -- CP-element group 260: 	167 
    -- CP-element group 260: 	171 
    -- CP-element group 260: 	159 
    -- CP-element group 260: 	163 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_Sample/ra
      -- 
    ra_8890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3510_inst_ack_0, ack => sendModule_CP_7961_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3510_Update/ca
      -- 
    ca_8895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3510_inst_ack_1, ack => sendModule_CP_7961_elements(261)); -- 
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	257 
    -- CP-element group 262: 	261 
    -- CP-element group 262: 	283 
    -- CP-element group 262: 	284 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	264 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (9) 
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/ptr_deref_3503_Split/$entry
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/ptr_deref_3503_Split/$exit
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/ptr_deref_3503_Split/split_req
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/ptr_deref_3503_Split/split_ack
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/word_access_start/$entry
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/word_access_start/word_0/$entry
      -- CP-element group 262: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/word_access_start/word_0/rr
      -- 
    rr_8933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(262), ack => ptr_deref_3503_store_0_req_0); -- 
    sendModule_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(257) & sendModule_CP_7961_elements(261) & sendModule_CP_7961_elements(283) & sendModule_CP_7961_elements(284) & sendModule_CP_7961_elements(264);
      gj_sendModule_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	265 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (5) 
      -- CP-element group 263: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_update_start_
      -- CP-element group 263: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Update/word_access_complete/$entry
      -- CP-element group 263: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Update/word_access_complete/word_0/$entry
      -- CP-element group 263: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Update/word_access_complete/word_0/cr
      -- 
    cr_8944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(263), ack => ptr_deref_3503_store_0_req_1); -- 
    sendModule_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(265);
      gj_sendModule_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	285 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	255 
    -- CP-element group 264: 	259 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (5) 
      -- CP-element group 264: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/word_access_start/$exit
      -- CP-element group 264: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/word_access_start/word_0/$exit
      -- CP-element group 264: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Sample/word_access_start/word_0/ra
      -- 
    ra_8934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3503_store_0_ack_0, ack => sendModule_CP_7961_elements(264)); -- 
    -- CP-element group 265:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	286 
    -- CP-element group 265: marked-successors 
    -- CP-element group 265: 	263 
    -- CP-element group 265:  members (5) 
      -- CP-element group 265: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Update/word_access_complete/$exit
      -- CP-element group 265: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Update/word_access_complete/word_0/$exit
      -- CP-element group 265: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_Update/word_access_complete/word_0/ca
      -- 
    ca_8945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3503_store_0_ack_1, ack => sendModule_CP_7961_elements(265)); -- 
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	141 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_Sample/req
      -- 
    req_8953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(266), ack => W_fetch_addr2_3332_delayed_8_0_3512_inst_req_0); -- 
    sendModule_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(141) & sendModule_CP_7961_elements(268);
      gj_sendModule_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	276 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_update_start_
      -- CP-element group 267: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_Update/req
      -- 
    req_8958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(267), ack => W_fetch_addr2_3332_delayed_8_0_3512_inst_req_1); -- 
    sendModule_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(276);
      gj_sendModule_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	136 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_Sample/ack
      -- 
    ack_8954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr2_3332_delayed_8_0_3512_inst_ack_0, ack => sendModule_CP_7961_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	274 
    -- CP-element group 269:  members (19) 
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_word_addrgen/root_register_ack
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_word_addrgen/root_register_req
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_word_addrgen/$exit
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_word_addrgen/$entry
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_plus_offset/sum_rename_ack
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_plus_offset/sum_rename_req
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/assign_stmt_3514_Update/ack
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_word_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_root_address_calculated
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_address_resized
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_addr_resize/$entry
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_addr_resize/$exit
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_addr_resize/base_resize_req
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_addr_resize/base_resize_ack
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_plus_offset/$entry
      -- CP-element group 269: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_base_plus_offset/$exit
      -- 
    ack_8959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr2_3332_delayed_8_0_3512_inst_ack_1, ack => sendModule_CP_7961_elements(269)); -- 
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	249 
    -- CP-element group 270: 	253 
    -- CP-element group 270: 	237 
    -- CP-element group 270: 	241 
    -- CP-element group 270: 	245 
    -- CP-element group 270: 	225 
    -- CP-element group 270: 	229 
    -- CP-element group 270: 	233 
    -- CP-element group 270: 	181 
    -- CP-element group 270: 	185 
    -- CP-element group 270: 	189 
    -- CP-element group 270: 	177 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_Sample/rr
      -- 
    rr_8967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(270), ack => CONCAT_u32_u64_3523_inst_req_0); -- 
    sendModule_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(249) & sendModule_CP_7961_elements(253) & sendModule_CP_7961_elements(237) & sendModule_CP_7961_elements(241) & sendModule_CP_7961_elements(245) & sendModule_CP_7961_elements(225) & sendModule_CP_7961_elements(229) & sendModule_CP_7961_elements(233) & sendModule_CP_7961_elements(181) & sendModule_CP_7961_elements(185) & sendModule_CP_7961_elements(189) & sendModule_CP_7961_elements(177) & sendModule_CP_7961_elements(272);
      gj_sendModule_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: marked-predecessors 
    -- CP-element group 271: 	276 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_update_start_
      -- CP-element group 271: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_Update/cr
      -- 
    cr_8972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(271), ack => CONCAT_u32_u64_3523_inst_req_1); -- 
    sendModule_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(276);
      gj_sendModule_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	251 
    -- CP-element group 272: 	235 
    -- CP-element group 272: 	239 
    -- CP-element group 272: 	243 
    -- CP-element group 272: 	247 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	223 
    -- CP-element group 272: 	227 
    -- CP-element group 272: 	231 
    -- CP-element group 272: 	183 
    -- CP-element group 272: 	187 
    -- CP-element group 272: 	175 
    -- CP-element group 272: 	179 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_Sample/ra
      -- 
    ra_8968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3523_inst_ack_0, ack => sendModule_CP_7961_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/CONCAT_u32_u64_3523_Update/ca
      -- 
    ca_8973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3523_inst_ack_1, ack => sendModule_CP_7961_elements(273)); -- 
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	269 
    -- CP-element group 274: 	273 
    -- CP-element group 274: 	285 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (9) 
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/word_access_start/word_0/rr
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/word_access_start/word_0/$entry
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/word_access_start/$entry
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/ptr_deref_3516_Split/split_ack
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/ptr_deref_3516_Split/split_req
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/ptr_deref_3516_Split/$exit
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/ptr_deref_3516_Split/$entry
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_sample_start_
      -- 
    rr_9011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(274), ack => ptr_deref_3516_store_0_req_0); -- 
    sendModule_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(269) & sendModule_CP_7961_elements(273) & sendModule_CP_7961_elements(285) & sendModule_CP_7961_elements(276);
      gj_sendModule_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	277 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (5) 
      -- CP-element group 275: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Update/word_access_complete/$entry
      -- CP-element group 275: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Update/word_access_complete/word_0/cr
      -- CP-element group 275: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Update/word_access_complete/word_0/$entry
      -- CP-element group 275: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_update_start_
      -- 
    cr_9022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(275), ack => ptr_deref_3516_store_0_req_1); -- 
    sendModule_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(277);
      gj_sendModule_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	286 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	142 
    -- CP-element group 276: 	267 
    -- CP-element group 276: 	271 
    -- CP-element group 276: 	274 
    -- CP-element group 276: 	146 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/word_access_start/word_0/ra
      -- CP-element group 276: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/word_access_start/word_0/$exit
      -- CP-element group 276: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/word_access_start/$exit
      -- CP-element group 276: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ring_reenable_memory_space_0
      -- CP-element group 276: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_sample_completed_
      -- 
    ra_9012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3516_store_0_ack_0, ack => sendModule_CP_7961_elements(276)); -- 
    -- CP-element group 277:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	286 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	275 
    -- CP-element group 277:  members (5) 
      -- CP-element group 277: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Update/word_access_complete/$exit
      -- CP-element group 277: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Update/word_access_complete/word_0/ca
      -- CP-element group 277: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_Update/word_access_complete/word_0/$exit
      -- CP-element group 277: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3516_update_completed_
      -- 
    ca_9023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3516_store_0_ack_1, ack => sendModule_CP_7961_elements(277)); -- 
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	15 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_Sample/rr
      -- CP-element group 278: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_Sample/$entry
      -- 
    rr_9031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(278), ack => SUB_u16_u16_3528_inst_req_0); -- 
    sendModule_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(15) & sendModule_CP_7961_elements(280);
      gj_sendModule_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_Update/cr
      -- CP-element group 279: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_update_start_
      -- 
    cr_9036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(279), ack => SUB_u16_u16_3528_inst_req_1); -- 
    sendModule_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_7961_elements(281);
      gj_sendModule_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	278 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_sample_completed_
      -- CP-element group 280: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_Sample/ra
      -- CP-element group 280: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_Sample/$exit
      -- 
    ra_9032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3528_inst_ack_0, ack => sendModule_CP_7961_elements(280)); -- 
    -- CP-element group 281:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	16 
    -- CP-element group 281: marked-successors 
    -- CP-element group 281: 	279 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_Update/ca
      -- CP-element group 281: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/SUB_u16_u16_3528_update_completed_
      -- 
    ca_9037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3528_inst_ack_1, ack => sendModule_CP_7961_elements(281)); -- 
    -- CP-element group 282:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	15 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	16 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group sendModule_CP_7961_elements(282) is a control-delay.
    cp_element_282_delay: control_delay_element  generic map(name => " 282_delay", delay_value => 1)  port map(req => sendModule_CP_7961_elements(15), ack => sendModule_CP_7961_elements(282), clk => clk, reset =>reset);
    -- CP-element group 283:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	144 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	262 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3335_ptr_deref_3503_delay
      -- 
    -- Element group sendModule_CP_7961_elements(283) is a control-delay.
    cp_element_283_delay: control_delay_element  generic map(name => " 283_delay", delay_value => 1)  port map(req => sendModule_CP_7961_elements(144), ack => sendModule_CP_7961_elements(283), clk => clk, reset =>reset);
    -- CP-element group 284:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	148 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	262 
    -- CP-element group 284:  members (1) 
      -- CP-element group 284: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3339_ptr_deref_3503_delay
      -- 
    -- Element group sendModule_CP_7961_elements(284) is a control-delay.
    cp_element_284_delay: control_delay_element  generic map(name => " 284_delay", delay_value => 1)  port map(req => sendModule_CP_7961_elements(148), ack => sendModule_CP_7961_elements(284), clk => clk, reset =>reset);
    -- CP-element group 285:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	264 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	274 
    -- CP-element group 285:  members (1) 
      -- CP-element group 285: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/ptr_deref_3503_ptr_deref_3516_delay
      -- 
    -- Element group sendModule_CP_7961_elements(285) is a control-delay.
    cp_element_285_delay: control_delay_element  generic map(name => " 285_delay", delay_value => 1)  port map(req => sendModule_CP_7961_elements(264), ack => sendModule_CP_7961_elements(285), clk => clk, reset =>reset);
    -- CP-element group 286:  join  transition  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	131 
    -- CP-element group 286: 	127 
    -- CP-element group 286: 	138 
    -- CP-element group 286: 	18 
    -- CP-element group 286: 	265 
    -- CP-element group 286: 	276 
    -- CP-element group 286: 	277 
    -- CP-element group 286: 	123 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	12 
    -- CP-element group 286:  members (1) 
      -- CP-element group 286: 	 branch_block_stmt_3181/do_while_stmt_3197/do_while_stmt_3197_loop_body/$exit
      -- 
    sendModule_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_7961_elements(131) & sendModule_CP_7961_elements(127) & sendModule_CP_7961_elements(138) & sendModule_CP_7961_elements(18) & sendModule_CP_7961_elements(265) & sendModule_CP_7961_elements(276) & sendModule_CP_7961_elements(277) & sendModule_CP_7961_elements(123);
      gj_sendModule_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_7961_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	11 
    -- CP-element group 287: successors 
    -- CP-element group 287:  members (2) 
      -- CP-element group 287: 	 branch_block_stmt_3181/do_while_stmt_3197/loop_exit/ack
      -- CP-element group 287: 	 branch_block_stmt_3181/do_while_stmt_3197/loop_exit/$exit
      -- 
    ack_9046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3197_branch_ack_0, ack => sendModule_CP_7961_elements(287)); -- 
    -- CP-element group 288:  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	11 
    -- CP-element group 288: successors 
    -- CP-element group 288:  members (2) 
      -- CP-element group 288: 	 branch_block_stmt_3181/do_while_stmt_3197/loop_taken/ack
      -- CP-element group 288: 	 branch_block_stmt_3181/do_while_stmt_3197/loop_taken/$exit
      -- 
    ack_9050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3197_branch_ack_1, ack => sendModule_CP_7961_elements(288)); -- 
    -- CP-element group 289:  transition  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	9 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	1 
    -- CP-element group 289:  members (1) 
      -- CP-element group 289: 	 branch_block_stmt_3181/do_while_stmt_3197/$exit
      -- 
    sendModule_CP_7961_elements(289) <= sendModule_CP_7961_elements(9);
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	1 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_sample_completed_
      -- CP-element group 290: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_update_start_
      -- CP-element group 290: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_Sample/$exit
      -- CP-element group 290: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_Sample/ack
      -- CP-element group 290: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_Update/req
      -- 
    ack_9063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3540_inst_ack_0, ack => sendModule_CP_7961_elements(290)); -- 
    req_9067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_7961_elements(290), ack => WPIPE_input_done_pipe_3540_inst_req_1); -- 
    -- CP-element group 291:  transition  place  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (8) 
      -- CP-element group 291: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_Update/$exit
      -- CP-element group 291: 	 $exit
      -- CP-element group 291: 	 branch_block_stmt_3181/$exit
      -- CP-element group 291: 	 branch_block_stmt_3181/branch_block_stmt_3181__exit__
      -- CP-element group 291: 	 branch_block_stmt_3181/assign_stmt_3542__exit__
      -- CP-element group 291: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_update_completed_
      -- CP-element group 291: 	 branch_block_stmt_3181/assign_stmt_3542/$exit
      -- CP-element group 291: 	 branch_block_stmt_3181/assign_stmt_3542/WPIPE_input_done_pipe_3540_Update/ack
      -- 
    ack_9068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3540_inst_ack_1, ack => sendModule_CP_7961_elements(291)); -- 
    sendModule_do_while_stmt_3197_terminator_9051: loop_terminator -- 
      generic map (name => " sendModule_do_while_stmt_3197_terminator_9051", max_iterations_in_flight =>15) 
      port map(loop_body_exit => sendModule_CP_7961_elements(12),loop_continue => sendModule_CP_7961_elements(288),loop_terminate => sendModule_CP_7961_elements(287),loop_back => sendModule_CP_7961_elements(10),loop_exit => sendModule_CP_7961_elements(9),clk => clk, reset => reset); -- 
    phi_stmt_3199_phi_seq_8083_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7961_elements(27);
      sendModule_CP_7961_elements(30)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7961_elements(30);
      sendModule_CP_7961_elements(31)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7961_elements(32);
      sendModule_CP_7961_elements(28) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7961_elements(25);
      sendModule_CP_7961_elements(34)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7961_elements(36);
      sendModule_CP_7961_elements(35)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7961_elements(37);
      sendModule_CP_7961_elements(26) <= phi_mux_reqs(1);
      phi_stmt_3199_phi_seq_8083 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3199_phi_seq_8083") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7961_elements(17), 
          phi_sample_ack => sendModule_CP_7961_elements(23), 
          phi_update_req => sendModule_CP_7961_elements(19), 
          phi_update_ack => sendModule_CP_7961_elements(24), 
          phi_mux_ack => sendModule_CP_7961_elements(29), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3204_phi_seq_8137_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7961_elements(46);
      sendModule_CP_7961_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7961_elements(53);
      sendModule_CP_7961_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7961_elements(54);
      sendModule_CP_7961_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7961_elements(44);
      sendModule_CP_7961_elements(55)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7961_elements(57);
      sendModule_CP_7961_elements(56)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7961_elements(58);
      sendModule_CP_7961_elements(45) <= phi_mux_reqs(1);
      phi_stmt_3204_phi_seq_8137 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3204_phi_seq_8137") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7961_elements(40), 
          phi_sample_ack => sendModule_CP_7961_elements(41), 
          phi_update_req => sendModule_CP_7961_elements(42), 
          phi_update_ack => sendModule_CP_7961_elements(43), 
          phi_mux_ack => sendModule_CP_7961_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3209_phi_seq_8181_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7961_elements(67);
      sendModule_CP_7961_elements(70)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7961_elements(70);
      sendModule_CP_7961_elements(71)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7961_elements(72);
      sendModule_CP_7961_elements(68) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7961_elements(65);
      sendModule_CP_7961_elements(74)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7961_elements(76);
      sendModule_CP_7961_elements(75)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7961_elements(77);
      sendModule_CP_7961_elements(66) <= phi_mux_reqs(1);
      phi_stmt_3209_phi_seq_8181 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3209_phi_seq_8181") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7961_elements(61), 
          phi_sample_ack => sendModule_CP_7961_elements(62), 
          phi_update_req => sendModule_CP_7961_elements(63), 
          phi_update_ack => sendModule_CP_7961_elements(64), 
          phi_mux_ack => sendModule_CP_7961_elements(69), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3214_phi_seq_8225_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7961_elements(86);
      sendModule_CP_7961_elements(89)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7961_elements(89);
      sendModule_CP_7961_elements(90)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7961_elements(91);
      sendModule_CP_7961_elements(87) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7961_elements(84);
      sendModule_CP_7961_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7961_elements(95);
      sendModule_CP_7961_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7961_elements(96);
      sendModule_CP_7961_elements(85) <= phi_mux_reqs(1);
      phi_stmt_3214_phi_seq_8225 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3214_phi_seq_8225") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7961_elements(80), 
          phi_sample_ack => sendModule_CP_7961_elements(81), 
          phi_update_req => sendModule_CP_7961_elements(82), 
          phi_update_ack => sendModule_CP_7961_elements(83), 
          phi_mux_ack => sendModule_CP_7961_elements(88), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3219_phi_seq_8269_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_7961_elements(105);
      sendModule_CP_7961_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_7961_elements(108);
      sendModule_CP_7961_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_7961_elements(110);
      sendModule_CP_7961_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_7961_elements(103);
      sendModule_CP_7961_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_7961_elements(114);
      sendModule_CP_7961_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_7961_elements(115);
      sendModule_CP_7961_elements(104) <= phi_mux_reqs(1);
      phi_stmt_3219_phi_seq_8269 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3219_phi_seq_8269") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_7961_elements(99), 
          phi_sample_ack => sendModule_CP_7961_elements(100), 
          phi_update_req => sendModule_CP_7961_elements(101), 
          phi_update_ack => sendModule_CP_7961_elements(102), 
          phi_mux_ack => sendModule_CP_7961_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_8035_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= sendModule_CP_7961_elements(13);
        preds(1)  <= sendModule_CP_7961_elements(14);
        entry_tmerge_8035 : transition_merge -- 
          generic map(name => " entry_tmerge_8035")
          port map (preds => preds, symbol_out => sendModule_CP_7961_elements(15));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_3247_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3256_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3265_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_3294_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3304_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3308_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3506_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3509_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3519_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3522_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_3510_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_3523_wire : std_logic_vector(63 downto 0);
    signal EQ_u2_u1_3261_3261_delayed_14_0_3391 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3269_3269_delayed_14_0_3405 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3277_3277_delayed_14_0_3419 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3285_3285_delayed_14_0_3433 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3293_3293_delayed_14_0_3447 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3301_3301_delayed_14_0_3461 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3309_3309_delayed_14_0_3475 : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_3317_3317_delayed_14_0_3489 : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_3318_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_3328_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_3194_wire : std_logic_vector(15 downto 0);
    signal MUX_3258_wire : std_logic_vector(15 downto 0);
    signal MUX_3296_wire : std_logic_vector(31 downto 0);
    signal MUX_3310_wire : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_3535_wire : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_3115_3115_delayed_1_0_3234 : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_3346_3346_delayed_1_0_3529 : std_logic_vector(15 downto 0);
    signal UGE_u16_u1_3239_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_3533_wire : std_logic_vector(0 downto 0);
    signal address1_3199 : std_logic_vector(31 downto 0);
    signal address2_3204 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3320_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3320_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3320_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3320_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3320_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3320_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3330_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3330_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3330_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3330_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3330_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3330_root_address : std_logic_vector(13 downto 0);
    signal cb_3187 : std_logic_vector(15 downto 0);
    signal chl_3209 : std_logic_vector(15 downto 0);
    signal chl_change_3241 : std_logic_vector(0 downto 0);
    signal chl_out_3190 : std_logic_vector(15 downto 0);
    signal col_3214 : std_logic_vector(15 downto 0);
    signal continue_flag_3537 : std_logic_vector(0 downto 0);
    signal fetch_addr1_3322 : std_logic_vector(31 downto 0);
    signal fetch_addr1_3322_delayed_8_0_3501 : std_logic_vector(31 downto 0);
    signal fetch_addr2_3332 : std_logic_vector(31 downto 0);
    signal fetch_addr2_3332_delayed_8_0_3514 : std_logic_vector(31 downto 0);
    signal fetch_val1_3336 : std_logic_vector(63 downto 0);
    signal fetch_val2_3340 : std_logic_vector(63 downto 0);
    signal konst_3232_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3244_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3246_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3252_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3255_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3264_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3317_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3327_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3389_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3403_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3417_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3431_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3445_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3459_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3473_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3487_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3527_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3541_wire_constant : std_logic_vector(7 downto 0);
    signal location1_3382 : std_logic_vector(1 downto 0);
    signal location2_3386 : std_logic_vector(1 downto 0);
    signal n_address1_3298 : std_logic_vector(31 downto 0);
    signal n_address1_3298_3203_buffered : std_logic_vector(31 downto 0);
    signal n_address2_3312 : std_logic_vector(31 downto 0);
    signal n_address2_3312_3208_buffered : std_logic_vector(31 downto 0);
    signal n_chl_3268 : std_logic_vector(15 downto 0);
    signal n_chl_3268_3213_buffered : std_logic_vector(15 downto 0);
    signal n_col_3249 : std_logic_vector(15 downto 0);
    signal n_col_3249_3218_buffered : std_logic_vector(15 downto 0);
    signal n_row_3260 : std_logic_vector(15 downto 0);
    signal n_row_3260_3223_buffered : std_logic_vector(15 downto 0);
    signal output_data1_3262_delayed_14_0_3394 : std_logic_vector(15 downto 0);
    signal output_data1_3270_delayed_14_0_3408 : std_logic_vector(15 downto 0);
    signal output_data1_3278_delayed_14_0_3422 : std_logic_vector(15 downto 0);
    signal output_data1_3286_delayed_14_0_3436 : std_logic_vector(15 downto 0);
    signal output_data1_3343 : std_logic_vector(15 downto 0);
    signal output_data2_3294_delayed_14_0_3450 : std_logic_vector(15 downto 0);
    signal output_data2_3302_delayed_14_0_3464 : std_logic_vector(15 downto 0);
    signal output_data2_3310_delayed_14_0_3478 : std_logic_vector(15 downto 0);
    signal output_data2_3318_delayed_14_0_3492 : std_logic_vector(15 downto 0);
    signal output_data2_3346 : std_logic_vector(15 downto 0);
    signal ptr_deref_3335_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3335_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3335_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3335_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3335_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3339_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3339_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3339_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3339_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3339_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3503_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3503_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3503_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3503_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3503_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3503_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3516_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3516_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3516_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3516_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3516_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3516_word_offset_0 : std_logic_vector(13 downto 0);
    signal rb_3184 : std_logic_vector(15 downto 0);
    signal row_3219 : std_logic_vector(15 downto 0);
    signal row_change_3229 : std_logic_vector(0 downto 0);
    signal row_size_3196 : std_logic_vector(31 downto 0);
    signal tmp1_3277 : std_logic_vector(31 downto 0);
    signal tmp2_3286 : std_logic_vector(31 downto 0);
    signal type_cast_3149_3149_delayed_1_0_3272 : std_logic_vector(31 downto 0);
    signal type_cast_3155_3155_delayed_1_0_3281 : std_logic_vector(31 downto 0);
    signal type_cast_3202_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3207_wire : std_logic_vector(31 downto 0);
    signal type_cast_3212_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3217_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3222_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3290_wire : std_logic_vector(31 downto 0);
    signal type_cast_3302_wire : std_logic_vector(31 downto 0);
    signal type_cast_3319_resized : std_logic_vector(13 downto 0);
    signal type_cast_3319_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3319_wire : std_logic_vector(63 downto 0);
    signal type_cast_3329_resized : std_logic_vector(13 downto 0);
    signal type_cast_3329_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3329_wire : std_logic_vector(63 downto 0);
    signal w11_3350 : std_logic_vector(15 downto 0);
    signal w12_3354 : std_logic_vector(15 downto 0);
    signal w13_3358 : std_logic_vector(15 downto 0);
    signal w14_3362 : std_logic_vector(15 downto 0);
    signal w21_3366 : std_logic_vector(15 downto 0);
    signal w22_3370 : std_logic_vector(15 downto 0);
    signal w23_3374 : std_logic_vector(15 downto 0);
    signal w24_3378 : std_logic_vector(15 downto 0);
    signal wb11_3400 : std_logic_vector(15 downto 0);
    signal wb12_3414 : std_logic_vector(15 downto 0);
    signal wb13_3428 : std_logic_vector(15 downto 0);
    signal wb14_3442 : std_logic_vector(15 downto 0);
    signal wb21_3456 : std_logic_vector(15 downto 0);
    signal wb22_3470 : std_logic_vector(15 downto 0);
    signal wb23_3484 : std_logic_vector(15 downto 0);
    signal wb24_3498 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_3320_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3320_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3320_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3320_resized_base_address <= "00000000000000";
    array_obj_ref_3330_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3330_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3330_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3330_resized_base_address <= "00000000000000";
    konst_3232_wire_constant <= "0000000000000001";
    konst_3244_wire_constant <= "0000000000000001";
    konst_3246_wire_constant <= "0000000000000001";
    konst_3252_wire_constant <= "0000000000000001";
    konst_3255_wire_constant <= "0000000000000010";
    konst_3264_wire_constant <= "0000000000000001";
    konst_3317_wire_constant <= "00000000000000000000000000000010";
    konst_3327_wire_constant <= "00000000000000000000000000000010";
    konst_3389_wire_constant <= "00";
    konst_3403_wire_constant <= "01";
    konst_3417_wire_constant <= "10";
    konst_3431_wire_constant <= "11";
    konst_3445_wire_constant <= "00";
    konst_3459_wire_constant <= "01";
    konst_3473_wire_constant <= "10";
    konst_3487_wire_constant <= "11";
    konst_3527_wire_constant <= "0000000000000001";
    konst_3541_wire_constant <= "00000001";
    ptr_deref_3335_word_offset_0 <= "00000000000000";
    ptr_deref_3339_word_offset_0 <= "00000000000000";
    ptr_deref_3503_word_offset_0 <= "00000000000000";
    ptr_deref_3516_word_offset_0 <= "00000000000000";
    type_cast_3202_wire_constant <= "00000000000000000000000000000000";
    type_cast_3212_wire_constant <= "0000000000000000";
    type_cast_3217_wire_constant <= "0000000000000001";
    type_cast_3222_wire_constant <= "0000000000000001";
    phi_stmt_3199: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3202_wire_constant & n_address1_3298_3203_buffered;
      req <= phi_stmt_3199_req_0 & phi_stmt_3199_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3199",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3199_ack_0,
          idata => idata,
          odata => address1_3199,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3199
    phi_stmt_3204: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3207_wire & n_address2_3312_3208_buffered;
      req <= phi_stmt_3204_req_0 & phi_stmt_3204_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3204",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3204_ack_0,
          idata => idata,
          odata => address2_3204,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3204
    phi_stmt_3209: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3212_wire_constant & n_chl_3268_3213_buffered;
      req <= phi_stmt_3209_req_0 & phi_stmt_3209_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3209",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3209_ack_0,
          idata => idata,
          odata => chl_3209,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3209
    phi_stmt_3214: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3217_wire_constant & n_col_3249_3218_buffered;
      req <= phi_stmt_3214_req_0 & phi_stmt_3214_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3214",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3214_ack_0,
          idata => idata,
          odata => col_3214,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3214
    phi_stmt_3219: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3222_wire_constant & n_row_3260_3223_buffered;
      req <= phi_stmt_3219_req_0 & phi_stmt_3219_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3219",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3219_ack_0,
          idata => idata,
          odata => row_3219,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3219
    -- flow-through select operator MUX_3248_inst
    n_col_3249 <= konst_3244_wire_constant when (row_change_3229(0) /=  '0') else ADD_u16_u16_3247_wire;
    -- flow-through select operator MUX_3258_inst
    MUX_3258_wire <= ADD_u16_u16_3256_wire when (row_change_3229(0) /=  '0') else row_3219;
    -- flow-through select operator MUX_3259_inst
    n_row_3260 <= konst_3252_wire_constant when (chl_change_3241(0) /=  '0') else MUX_3258_wire;
    -- flow-through select operator MUX_3267_inst
    n_chl_3268 <= ADD_u16_u16_3265_wire when (chl_change_3241(0) /=  '0') else chl_3209;
    -- flow-through select operator MUX_3296_inst
    MUX_3296_wire <= ADD_u32_u32_3294_wire when (row_change_3229(0) /=  '0') else tmp1_3277;
    -- flow-through select operator MUX_3297_inst
    n_address1_3298 <= type_cast_3290_wire when (chl_change_3241(0) /=  '0') else MUX_3296_wire;
    -- flow-through select operator MUX_3310_inst
    MUX_3310_wire <= ADD_u32_u32_3308_wire when (row_change_3229(0) /=  '0') else tmp2_3286;
    -- flow-through select operator MUX_3311_inst
    n_address2_3312 <= ADD_u32_u32_3304_wire when (chl_change_3241(0) /=  '0') else MUX_3310_wire;
    -- flow-through select operator MUX_3399_inst
    wb11_3400 <= output_data1_3262_delayed_14_0_3394 when (EQ_u2_u1_3261_3261_delayed_14_0_3391(0) /=  '0') else w11_3350;
    -- flow-through select operator MUX_3413_inst
    wb12_3414 <= output_data1_3270_delayed_14_0_3408 when (EQ_u2_u1_3269_3269_delayed_14_0_3405(0) /=  '0') else w12_3354;
    -- flow-through select operator MUX_3427_inst
    wb13_3428 <= output_data1_3278_delayed_14_0_3422 when (EQ_u2_u1_3277_3277_delayed_14_0_3419(0) /=  '0') else w13_3358;
    -- flow-through select operator MUX_3441_inst
    wb14_3442 <= output_data1_3286_delayed_14_0_3436 when (EQ_u2_u1_3285_3285_delayed_14_0_3433(0) /=  '0') else w14_3362;
    -- flow-through select operator MUX_3455_inst
    wb21_3456 <= output_data2_3294_delayed_14_0_3450 when (EQ_u2_u1_3293_3293_delayed_14_0_3447(0) /=  '0') else w21_3366;
    -- flow-through select operator MUX_3469_inst
    wb22_3470 <= output_data2_3302_delayed_14_0_3464 when (EQ_u2_u1_3301_3301_delayed_14_0_3461(0) /=  '0') else w22_3370;
    -- flow-through select operator MUX_3483_inst
    wb23_3484 <= output_data2_3310_delayed_14_0_3478 when (EQ_u2_u1_3309_3309_delayed_14_0_3475(0) /=  '0') else w23_3374;
    -- flow-through select operator MUX_3497_inst
    wb24_3498 <= output_data2_3318_delayed_14_0_3492 when (EQ_u2_u1_3317_3317_delayed_14_0_3489(0) /=  '0') else w24_3378;
    slice_3349_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3349_inst_req_0;
      slice_3349_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3349_inst_req_1;
      slice_3349_inst_ack_1<= update_ack(0);
      slice_3349_inst: SliceSplitProtocol generic map(name => "slice_3349_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3336, dout => w11_3350, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3353_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3353_inst_req_0;
      slice_3353_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3353_inst_req_1;
      slice_3353_inst_ack_1<= update_ack(0);
      slice_3353_inst: SliceSplitProtocol generic map(name => "slice_3353_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3336, dout => w12_3354, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3357_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3357_inst_req_0;
      slice_3357_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3357_inst_req_1;
      slice_3357_inst_ack_1<= update_ack(0);
      slice_3357_inst: SliceSplitProtocol generic map(name => "slice_3357_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3336, dout => w13_3358, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3361_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3361_inst_req_0;
      slice_3361_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3361_inst_req_1;
      slice_3361_inst_ack_1<= update_ack(0);
      slice_3361_inst: SliceSplitProtocol generic map(name => "slice_3361_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3336, dout => w14_3362, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3365_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3365_inst_req_0;
      slice_3365_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3365_inst_req_1;
      slice_3365_inst_ack_1<= update_ack(0);
      slice_3365_inst: SliceSplitProtocol generic map(name => "slice_3365_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3340, dout => w21_3366, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3369_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3369_inst_req_0;
      slice_3369_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3369_inst_req_1;
      slice_3369_inst_ack_1<= update_ack(0);
      slice_3369_inst: SliceSplitProtocol generic map(name => "slice_3369_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3340, dout => w22_3370, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3373_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3373_inst_req_0;
      slice_3373_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3373_inst_req_1;
      slice_3373_inst_ack_1<= update_ack(0);
      slice_3373_inst: SliceSplitProtocol generic map(name => "slice_3373_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3340, dout => w23_3374, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3377_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3377_inst_req_0;
      slice_3377_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3377_inst_req_1;
      slice_3377_inst_ack_1<= update_ack(0);
      slice_3377_inst: SliceSplitProtocol generic map(name => "slice_3377_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3340, dout => w24_3378, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_fetch_addr1_3322_delayed_8_0_3499_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr1_3322_delayed_8_0_3499_inst_req_0;
      W_fetch_addr1_3322_delayed_8_0_3499_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr1_3322_delayed_8_0_3499_inst_req_1;
      W_fetch_addr1_3322_delayed_8_0_3499_inst_ack_1<= rack(0);
      W_fetch_addr1_3322_delayed_8_0_3499_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr1_3322_delayed_8_0_3499_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr1_3322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_3322_delayed_8_0_3501,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_addr2_3332_delayed_8_0_3512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr2_3332_delayed_8_0_3512_inst_req_0;
      W_fetch_addr2_3332_delayed_8_0_3512_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr2_3332_delayed_8_0_3512_inst_req_1;
      W_fetch_addr2_3332_delayed_8_0_3512_inst_ack_1<= rack(0);
      W_fetch_addr2_3332_delayed_8_0_3512_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr2_3332_delayed_8_0_3512_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr2_3332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_3332_delayed_8_0_3514,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3262_delayed_14_0_3392_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3262_delayed_14_0_3392_inst_req_0;
      W_output_data1_3262_delayed_14_0_3392_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3262_delayed_14_0_3392_inst_req_1;
      W_output_data1_3262_delayed_14_0_3392_inst_ack_1<= rack(0);
      W_output_data1_3262_delayed_14_0_3392_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3262_delayed_14_0_3392_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3262_delayed_14_0_3394,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3270_delayed_14_0_3406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3270_delayed_14_0_3406_inst_req_0;
      W_output_data1_3270_delayed_14_0_3406_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3270_delayed_14_0_3406_inst_req_1;
      W_output_data1_3270_delayed_14_0_3406_inst_ack_1<= rack(0);
      W_output_data1_3270_delayed_14_0_3406_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3270_delayed_14_0_3406_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3270_delayed_14_0_3408,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3278_delayed_14_0_3420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3278_delayed_14_0_3420_inst_req_0;
      W_output_data1_3278_delayed_14_0_3420_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3278_delayed_14_0_3420_inst_req_1;
      W_output_data1_3278_delayed_14_0_3420_inst_ack_1<= rack(0);
      W_output_data1_3278_delayed_14_0_3420_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3278_delayed_14_0_3420_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3278_delayed_14_0_3422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3286_delayed_14_0_3434_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3286_delayed_14_0_3434_inst_req_0;
      W_output_data1_3286_delayed_14_0_3434_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3286_delayed_14_0_3434_inst_req_1;
      W_output_data1_3286_delayed_14_0_3434_inst_ack_1<= rack(0);
      W_output_data1_3286_delayed_14_0_3434_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3286_delayed_14_0_3434_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3286_delayed_14_0_3436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3294_delayed_14_0_3448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3294_delayed_14_0_3448_inst_req_0;
      W_output_data2_3294_delayed_14_0_3448_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3294_delayed_14_0_3448_inst_req_1;
      W_output_data2_3294_delayed_14_0_3448_inst_ack_1<= rack(0);
      W_output_data2_3294_delayed_14_0_3448_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3294_delayed_14_0_3448_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3294_delayed_14_0_3450,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3302_delayed_14_0_3462_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3302_delayed_14_0_3462_inst_req_0;
      W_output_data2_3302_delayed_14_0_3462_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3302_delayed_14_0_3462_inst_req_1;
      W_output_data2_3302_delayed_14_0_3462_inst_ack_1<= rack(0);
      W_output_data2_3302_delayed_14_0_3462_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3302_delayed_14_0_3462_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3302_delayed_14_0_3464,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3310_delayed_14_0_3476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3310_delayed_14_0_3476_inst_req_0;
      W_output_data2_3310_delayed_14_0_3476_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3310_delayed_14_0_3476_inst_req_1;
      W_output_data2_3310_delayed_14_0_3476_inst_ack_1<= rack(0);
      W_output_data2_3310_delayed_14_0_3476_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3310_delayed_14_0_3476_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3310_delayed_14_0_3478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3318_delayed_14_0_3490_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3318_delayed_14_0_3490_inst_req_0;
      W_output_data2_3318_delayed_14_0_3490_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3318_delayed_14_0_3490_inst_req_1;
      W_output_data2_3318_delayed_14_0_3490_inst_ack_1<= rack(0);
      W_output_data2_3318_delayed_14_0_3490_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3318_delayed_14_0_3490_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3318_delayed_14_0_3492,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3321_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3321_final_reg_req_0;
      addr_of_3321_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3321_final_reg_req_1;
      addr_of_3321_final_reg_ack_1<= rack(0);
      addr_of_3321_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3321_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3320_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_3322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3331_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3331_final_reg_req_0;
      addr_of_3331_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3331_final_reg_req_1;
      addr_of_3331_final_reg_ack_1<= rack(0);
      addr_of_3331_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3331_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3330_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_3332,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_3298_3203_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_3298_3203_buf_req_0;
      n_address1_3298_3203_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_3298_3203_buf_req_1;
      n_address1_3298_3203_buf_ack_1<= rack(0);
      n_address1_3298_3203_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_3298_3203_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_3298,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_3298_3203_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_3312_3208_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_3312_3208_buf_req_0;
      n_address2_3312_3208_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_3312_3208_buf_req_1;
      n_address2_3312_3208_buf_ack_1<= rack(0);
      n_address2_3312_3208_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_3312_3208_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_3312,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_3312_3208_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_3268_3213_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_3268_3213_buf_req_0;
      n_chl_3268_3213_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_3268_3213_buf_req_1;
      n_chl_3268_3213_buf_ack_1<= rack(0);
      n_chl_3268_3213_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_3268_3213_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_3268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_3268_3213_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_3249_3218_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_3249_3218_buf_req_0;
      n_col_3249_3218_buf_ack_0<= wack(0);
      rreq(0) <= n_col_3249_3218_buf_req_1;
      n_col_3249_3218_buf_ack_1<= rack(0);
      n_col_3249_3218_buf : InterlockBuffer generic map ( -- 
        name => "n_col_3249_3218_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_3249,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_3249_3218_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_3260_3223_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_3260_3223_buf_req_0;
      n_row_3260_3223_buf_ack_0<= wack(0);
      rreq(0) <= n_row_3260_3223_buf_req_1;
      n_row_3260_3223_buf_ack_1<= rack(0);
      n_row_3260_3223_buf : InterlockBuffer generic map ( -- 
        name => "n_row_3260_3223_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_3260,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_3260_3223_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3195_inst
    process(MUL_u16_u16_3194_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_3194_wire(15 downto 0);
      row_size_3196 <= tmp_var; -- 
    end process;
    type_cast_3207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3207_inst_req_0;
      type_cast_3207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3207_inst_req_1;
      type_cast_3207_inst_ack_1<= rack(0);
      type_cast_3207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => row_size_3196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3207_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3271_inst_req_0;
      type_cast_3271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3271_inst_req_1;
      type_cast_3271_inst_ack_1<= rack(0);
      type_cast_3271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3271_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_3190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3149_3149_delayed_1_0_3272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3280_inst_req_0;
      type_cast_3280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3280_inst_req_1;
      type_cast_3280_inst_ack_1<= rack(0);
      type_cast_3280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3280_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_3190,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3155_3155_delayed_1_0_3281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3290_inst
    process(n_chl_3268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3268(15 downto 0);
      type_cast_3290_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3302_inst
    process(n_chl_3268) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3268(15 downto 0);
      type_cast_3302_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3319_inst
    process(LSHR_u32_u32_3318_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3318_wire(31 downto 0);
      type_cast_3319_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3329_inst
    process(LSHR_u32_u32_3328_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3328_wire(31 downto 0);
      type_cast_3329_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3381_inst
    process(address1_3199) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := address1_3199(1 downto 0);
      location1_3382 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3385_inst
    process(address2_3204) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := address2_3204(1 downto 0);
      location2_3386 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_3320_index_1_rename
    process(type_cast_3319_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3319_resized;
      ov(13 downto 0) := iv;
      type_cast_3319_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3320_index_1_resize
    process(type_cast_3319_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3319_wire;
      ov := iv(13 downto 0);
      type_cast_3319_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3320_root_address_inst
    process(array_obj_ref_3320_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3320_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3320_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3330_index_1_rename
    process(type_cast_3329_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3329_resized;
      ov(13 downto 0) := iv;
      type_cast_3329_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3330_index_1_resize
    process(type_cast_3329_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3329_wire;
      ov := iv(13 downto 0);
      type_cast_3329_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3330_root_address_inst
    process(array_obj_ref_3330_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3330_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3330_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3335_addr_0
    process(ptr_deref_3335_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3335_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3335_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3335_base_resize
    process(fetch_addr1_3322) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_3322;
      ov := iv(13 downto 0);
      ptr_deref_3335_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3335_gather_scatter
    process(ptr_deref_3335_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3335_data_0;
      ov(63 downto 0) := iv;
      fetch_val1_3336 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3335_root_address_inst
    process(ptr_deref_3335_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3335_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3335_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3339_addr_0
    process(ptr_deref_3339_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3339_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3339_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3339_base_resize
    process(fetch_addr2_3332) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_3332;
      ov := iv(13 downto 0);
      ptr_deref_3339_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3339_gather_scatter
    process(ptr_deref_3339_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3339_data_0;
      ov(63 downto 0) := iv;
      fetch_val2_3340 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3339_root_address_inst
    process(ptr_deref_3339_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3339_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3339_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3503_addr_0
    process(ptr_deref_3503_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3503_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3503_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3503_base_resize
    process(fetch_addr1_3322_delayed_8_0_3501) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_3322_delayed_8_0_3501;
      ov := iv(13 downto 0);
      ptr_deref_3503_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3503_gather_scatter
    process(CONCAT_u32_u64_3510_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3510_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3503_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3503_root_address_inst
    process(ptr_deref_3503_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3503_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3503_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3516_addr_0
    process(ptr_deref_3516_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3516_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3516_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3516_base_resize
    process(fetch_addr2_3332_delayed_8_0_3514) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_3332_delayed_8_0_3514;
      ov := iv(13 downto 0);
      ptr_deref_3516_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3516_gather_scatter
    process(CONCAT_u32_u64_3523_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3523_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3516_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3516_root_address_inst
    process(ptr_deref_3516_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3516_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3516_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_3197_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_3537;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3197_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3197_branch_req_0,
          ack0 => do_while_stmt_3197_branch_ack_0,
          ack1 => do_while_stmt_3197_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3247_inst
    process(col_3214) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_3214, konst_3246_wire_constant, tmp_var);
      ADD_u16_u16_3247_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3256_inst
    process(row_3219) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_3219, konst_3255_wire_constant, tmp_var);
      ADD_u16_u16_3256_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3265_inst
    process(chl_3209) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_3209, konst_3264_wire_constant, tmp_var);
      ADD_u16_u16_3265_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3276_inst
    process(address1_3199, type_cast_3149_3149_delayed_1_0_3272) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_3199, type_cast_3149_3149_delayed_1_0_3272, tmp_var);
      tmp1_3277 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3285_inst
    process(address2_3204, type_cast_3155_3155_delayed_1_0_3281) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_3204, type_cast_3155_3155_delayed_1_0_3281, tmp_var);
      tmp2_3286 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3294_inst
    process(tmp1_3277, row_size_3196) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_3277, row_size_3196, tmp_var);
      ADD_u32_u32_3294_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3304_inst
    process(type_cast_3302_wire, row_size_3196) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_3302_wire, row_size_3196, tmp_var);
      ADD_u32_u32_3304_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3308_inst
    process(tmp2_3286, row_size_3196) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_3286, row_size_3196, tmp_var);
      ADD_u32_u32_3308_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3240_inst
    process(row_change_3229, UGE_u16_u1_3239_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(row_change_3229, UGE_u16_u1_3239_wire, tmp_var);
      chl_change_3241 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3506_inst
    process(wb11_3400, wb12_3414) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb11_3400, wb12_3414, tmp_var);
      CONCAT_u16_u32_3506_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3509_inst
    process(wb13_3428, wb14_3442) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb13_3428, wb14_3442, tmp_var);
      CONCAT_u16_u32_3509_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3519_inst
    process(wb21_3456, wb22_3470) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb21_3456, wb22_3470, tmp_var);
      CONCAT_u16_u32_3519_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3522_inst
    process(wb23_3484, wb24_3498) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(wb23_3484, wb24_3498, tmp_var);
      CONCAT_u16_u32_3522_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : CONCAT_u32_u64_3510_inst 
    ApConcat_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3506_wire & CONCAT_u16_u32_3509_wire;
      CONCAT_u32_u64_3510_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3510_inst_req_0;
      CONCAT_u32_u64_3510_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3510_inst_req_1;
      CONCAT_u32_u64_3510_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_13_gI: SplitGuardInterface generic map(name => "ApConcat_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : CONCAT_u32_u64_3523_inst 
    ApConcat_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3519_wire & CONCAT_u16_u32_3522_wire;
      CONCAT_u32_u64_3523_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3523_inst_req_0;
      CONCAT_u32_u64_3523_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3523_inst_req_1;
      CONCAT_u32_u64_3523_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_14_gI: SplitGuardInterface generic map(name => "ApConcat_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- binary operator EQ_u16_u1_3228_inst
    process(col_3214, cb_3187) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_3214, cb_3187, tmp_var);
      row_change_3229 <= tmp_var; --
    end process;
    -- shared split operator group (16) : EQ_u2_u1_3390_inst 
    ApIntEq_group_16: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3382;
      EQ_u2_u1_3261_3261_delayed_14_0_3391 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3390_inst_req_0;
      EQ_u2_u1_3390_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3390_inst_req_1;
      EQ_u2_u1_3390_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_16_gI: SplitGuardInterface generic map(name => "ApIntEq_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : EQ_u2_u1_3404_inst 
    ApIntEq_group_17: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3382;
      EQ_u2_u1_3269_3269_delayed_14_0_3405 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3404_inst_req_0;
      EQ_u2_u1_3404_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3404_inst_req_1;
      EQ_u2_u1_3404_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_17_gI: SplitGuardInterface generic map(name => "ApIntEq_group_17_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_17",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : EQ_u2_u1_3418_inst 
    ApIntEq_group_18: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3382;
      EQ_u2_u1_3277_3277_delayed_14_0_3419 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3418_inst_req_0;
      EQ_u2_u1_3418_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3418_inst_req_1;
      EQ_u2_u1_3418_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_18_gI: SplitGuardInterface generic map(name => "ApIntEq_group_18_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_18",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "10",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : EQ_u2_u1_3432_inst 
    ApIntEq_group_19: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3382;
      EQ_u2_u1_3285_3285_delayed_14_0_3433 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3432_inst_req_0;
      EQ_u2_u1_3432_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3432_inst_req_1;
      EQ_u2_u1_3432_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_19_gI: SplitGuardInterface generic map(name => "ApIntEq_group_19_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_19",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : EQ_u2_u1_3446_inst 
    ApIntEq_group_20: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3386;
      EQ_u2_u1_3293_3293_delayed_14_0_3447 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3446_inst_req_0;
      EQ_u2_u1_3446_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3446_inst_req_1;
      EQ_u2_u1_3446_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_20_gI: SplitGuardInterface generic map(name => "ApIntEq_group_20_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_20",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : EQ_u2_u1_3460_inst 
    ApIntEq_group_21: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3386;
      EQ_u2_u1_3301_3301_delayed_14_0_3461 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3460_inst_req_0;
      EQ_u2_u1_3460_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3460_inst_req_1;
      EQ_u2_u1_3460_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_21_gI: SplitGuardInterface generic map(name => "ApIntEq_group_21_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_21",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : EQ_u2_u1_3474_inst 
    ApIntEq_group_22: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3386;
      EQ_u2_u1_3309_3309_delayed_14_0_3475 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3474_inst_req_0;
      EQ_u2_u1_3474_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3474_inst_req_1;
      EQ_u2_u1_3474_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_22_gI: SplitGuardInterface generic map(name => "ApIntEq_group_22_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_22",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "10",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : EQ_u2_u1_3488_inst 
    ApIntEq_group_23: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3386;
      EQ_u2_u1_3317_3317_delayed_14_0_3489 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u2_u1_3488_inst_req_0;
      EQ_u2_u1_3488_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u2_u1_3488_inst_req_1;
      EQ_u2_u1_3488_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_23_gI: SplitGuardInterface generic map(name => "ApIntEq_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 2,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11",
          constant_width => 2,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- binary operator LSHR_u32_u32_3318_inst
    process(address1_3199) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_3199, konst_3317_wire_constant, tmp_var);
      LSHR_u32_u32_3318_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3328_inst
    process(address2_3204) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_3204, konst_3327_wire_constant, tmp_var);
      LSHR_u32_u32_3328_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3194_inst
    process(chl_out_3190, cb_3187) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_out_3190, cb_3187, tmp_var);
      MUL_u16_u16_3194_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_3535_inst
    process(chl_change_3241) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", chl_change_3241, tmp_var);
      NOT_u1_u1_3535_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_3536_inst
    process(ULT_u16_u1_3533_wire, NOT_u1_u1_3535_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ULT_u16_u1_3533_wire, NOT_u1_u1_3535_wire, tmp_var);
      continue_flag_3537 <= tmp_var; --
    end process;
    -- shared split operator group (29) : SUB_u16_u16_3233_inst 
    ApIntSub_group_29: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rb_3184;
      SUB_u16_u16_3115_3115_delayed_1_0_3234 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3233_inst_req_0;
      SUB_u16_u16_3233_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3233_inst_req_1;
      SUB_u16_u16_3233_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_29_gI: SplitGuardInterface generic map(name => "ApIntSub_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : SUB_u16_u16_3528_inst 
    ApIntSub_group_30: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= chl_out_3190;
      SUB_u16_u16_3346_3346_delayed_1_0_3529 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3528_inst_req_0;
      SUB_u16_u16_3528_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3528_inst_req_1;
      SUB_u16_u16_3528_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_30_gI: SplitGuardInterface generic map(name => "ApIntSub_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- binary operator UGE_u16_u1_3239_inst
    process(row_3219, SUB_u16_u16_3115_3115_delayed_1_0_3234) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(row_3219, SUB_u16_u16_3115_3115_delayed_1_0_3234, tmp_var);
      UGE_u16_u1_3239_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_3533_inst
    process(chl_3209, SUB_u16_u16_3346_3346_delayed_1_0_3529) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(chl_3209, SUB_u16_u16_3346_3346_delayed_1_0_3529, tmp_var);
      ULT_u16_u1_3533_wire <= tmp_var; --
    end process;
    -- shared split operator group (33) : array_obj_ref_3320_index_offset 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3319_scaled;
      array_obj_ref_3320_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3320_index_offset_req_0;
      array_obj_ref_3320_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3320_index_offset_req_1;
      array_obj_ref_3320_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : array_obj_ref_3330_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3329_scaled;
      array_obj_ref_3330_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3330_index_offset_req_0;
      array_obj_ref_3330_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3330_index_offset_req_1;
      array_obj_ref_3330_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared load operator group (0) : ptr_deref_3335_load_0 ptr_deref_3339_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3335_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3339_load_0_req_0;
      ptr_deref_3335_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3339_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3335_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3339_load_0_req_1;
      ptr_deref_3335_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3339_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3335_word_address_0 & ptr_deref_3339_word_address_0;
      ptr_deref_3335_data_0 <= data_out(127 downto 64);
      ptr_deref_3339_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3503_store_0 ptr_deref_3516_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3503_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3516_store_0_req_0;
      ptr_deref_3503_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3516_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3503_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3516_store_0_req_1;
      ptr_deref_3503_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3516_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3503_word_address_0 & ptr_deref_3516_word_address_0;
      data_in <= ptr_deref_3503_data_0 & ptr_deref_3516_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_output_pipe_3189_inst RPIPE_output_pipe_3186_inst RPIPE_output_pipe_3183_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(47 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 2 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= RPIPE_output_pipe_3189_inst_req_0;
      reqL_unguarded(1) <= RPIPE_output_pipe_3186_inst_req_0;
      reqL_unguarded(0) <= RPIPE_output_pipe_3183_inst_req_0;
      RPIPE_output_pipe_3189_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_output_pipe_3186_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_output_pipe_3183_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= RPIPE_output_pipe_3189_inst_req_1;
      reqR_unguarded(1) <= RPIPE_output_pipe_3186_inst_req_1;
      reqR_unguarded(0) <= RPIPE_output_pipe_3183_inst_req_1;
      RPIPE_output_pipe_3189_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_output_pipe_3186_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_output_pipe_3183_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      chl_out_3190 <= data_out(47 downto 32);
      cb_3187 <= data_out(31 downto 16);
      rb_3184 <= data_out(15 downto 0);
      output_pipe_read_0_gI: SplitGuardInterface generic map(name => "output_pipe_read_0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_0: InputPortRevised -- 
        generic map ( name => "output_pipe_read_0", data_width => 16,  num_reqs => 3,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(1),
          oack => output_pipe_pipe_read_ack(1),
          odata => output_pipe_pipe_read_data(31 downto 16),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_output_pipe_3342_inst RPIPE_output_pipe_3345_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_output_pipe_3342_inst_req_0;
      reqL_unguarded(0) <= RPIPE_output_pipe_3345_inst_req_0;
      RPIPE_output_pipe_3342_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_output_pipe_3345_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_output_pipe_3342_inst_req_1;
      reqR_unguarded(0) <= RPIPE_output_pipe_3345_inst_req_1;
      RPIPE_output_pipe_3342_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_output_pipe_3345_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      output_data1_3343 <= data_out(31 downto 16);
      output_data2_3346 <= data_out(15 downto 0);
      output_pipe_read_1_gI: SplitGuardInterface generic map(name => "output_pipe_read_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_1: InputPortRevised -- 
        generic map ( name => "output_pipe_read_1", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(0),
          oack => output_pipe_pipe_read_ack(0),
          odata => output_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3540_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3540_inst_req_0;
      WPIPE_input_done_pipe_3540_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3540_inst_req_1;
      WPIPE_input_done_pipe_3540_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3541_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendModule_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_1601_start: Boolean;
  signal timer_CP_1601_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_515_inst_ack_1 : boolean;
  signal WPIPE_timer_req_515_inst_req_1 : boolean;
  signal WPIPE_timer_req_515_inst_ack_0 : boolean;
  signal WPIPE_timer_req_515_inst_req_0 : boolean;
  signal RPIPE_timer_resp_520_inst_req_0 : boolean;
  signal RPIPE_timer_resp_520_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_520_inst_req_1 : boolean;
  signal RPIPE_timer_resp_520_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_1601_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1601_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_1601_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1601_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_1601: Block -- control-path 
    signal timer_CP_1601_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_1601_elements(0) <= timer_CP_1601_start;
    timer_CP_1601_symbol <= timer_CP_1601_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/$entry
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_sample_start_
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Sample/req
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_sample_start_
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Sample/rr
      -- 
    rr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1601_elements(0), ack => RPIPE_timer_resp_520_inst_req_0); -- 
    req_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1601_elements(0), ack => WPIPE_timer_req_515_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Update/req
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_sample_completed_
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Update/$entry
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Sample/ack
      -- CP-element group 1: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_update_start_
      -- 
    ack_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_515_inst_ack_0, ack => timer_CP_1601_elements(1)); -- 
    req_1619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1601_elements(1), ack => WPIPE_timer_req_515_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Update/ack
      -- CP-element group 2: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_Update/$exit
      -- CP-element group 2: 	 assign_stmt_518_to_assign_stmt_521/WPIPE_timer_req_515_update_completed_
      -- 
    ack_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_515_inst_ack_1, ack => timer_CP_1601_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_update_start_
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_sample_completed_
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Sample/ra
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Update/$entry
      -- CP-element group 3: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Update/cr
      -- 
    ra_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_520_inst_ack_0, ack => timer_CP_1601_elements(3)); -- 
    cr_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1601_elements(3), ack => RPIPE_timer_resp_520_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_update_completed_
      -- CP-element group 4: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Update/$exit
      -- CP-element group 4: 	 assign_stmt_518_to_assign_stmt_521/RPIPE_timer_resp_520_Update/ca
      -- 
    ca_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_520_inst_ack_1, ack => timer_CP_1601_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_518_to_assign_stmt_521/$exit
      -- CP-element group 5: 	 $exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_1601_elements(2) & timer_CP_1601_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_1601_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_517_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_517_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_520_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_520_inst_req_0;
      RPIPE_timer_resp_520_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_520_inst_req_1;
      RPIPE_timer_resp_520_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_515_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_515_inst_req_0;
      WPIPE_timer_req_515_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_515_inst_req_1;
      WPIPE_timer_req_515_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_517_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_9964_start: Boolean;
  signal timerDaemon_CP_9964_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nCOUNTER_3833_3824_buf_ack_0 : boolean;
  signal nCOUNTER_3833_3824_buf_req_0 : boolean;
  signal phi_stmt_3820_req_1 : boolean;
  signal WPIPE_timer_resp_3835_inst_req_1 : boolean;
  signal WPIPE_timer_resp_3835_inst_ack_1 : boolean;
  signal do_while_stmt_3818_branch_req_0 : boolean;
  signal phi_stmt_3820_ack_0 : boolean;
  signal phi_stmt_3820_req_0 : boolean;
  signal RPIPE_timer_req_3827_inst_req_0 : boolean;
  signal RPIPE_timer_req_3827_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_3835_inst_req_0 : boolean;
  signal WPIPE_timer_resp_3835_inst_ack_0 : boolean;
  signal nCOUNTER_3833_3824_buf_req_1 : boolean;
  signal nCOUNTER_3833_3824_buf_ack_1 : boolean;
  signal do_while_stmt_3818_branch_ack_1 : boolean;
  signal do_while_stmt_3818_branch_ack_0 : boolean;
  signal RPIPE_timer_req_3827_inst_req_1 : boolean;
  signal RPIPE_timer_req_3827_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_9964_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_9964_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_9964_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_9964_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_9964: Block -- control-path 
    signal timerDaemon_CP_9964_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_9964_elements(0) <= timerDaemon_CP_9964_start;
    timerDaemon_CP_9964_symbol <= timerDaemon_CP_9964_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_3817/do_while_stmt_3818__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3817/$entry
      -- CP-element group 0: 	 branch_block_stmt_3817/branch_block_stmt_3817__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_3817/do_while_stmt_3818__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_3817/$exit
      -- CP-element group 1: 	 branch_block_stmt_3817/branch_block_stmt_3817__exit__
      -- 
    timerDaemon_CP_9964_elements(1) <= timerDaemon_CP_9964_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_3817/do_while_stmt_3818/$entry
      -- CP-element group 2: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818__entry__
      -- 
    timerDaemon_CP_9964_elements(2) <= timerDaemon_CP_9964_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818__exit__
      -- 
    -- Element group timerDaemon_CP_9964_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_3817/do_while_stmt_3818/loop_back
      -- 
    -- Element group timerDaemon_CP_9964_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_3817/do_while_stmt_3818/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_3817/do_while_stmt_3818/condition_done
      -- CP-element group 5: 	 branch_block_stmt_3817/do_while_stmt_3818/loop_exit/$entry
      -- 
    timerDaemon_CP_9964_elements(5) <= timerDaemon_CP_9964_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_3817/do_while_stmt_3818/loop_body_done
      -- 
    timerDaemon_CP_9964_elements(6) <= timerDaemon_CP_9964_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_9964_elements(7) <= timerDaemon_CP_9964_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_9964_elements(8) <= timerDaemon_CP_9964_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3825_sample_start_
      -- 
    -- Element group timerDaemon_CP_9964_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/condition_evaluated
      -- 
    condition_evaluated_9988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_9988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(10), ack => do_while_stmt_3818_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(40) & timerDaemon_CP_9964_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/aggregated_phi_sample_req
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(9) & timerDaemon_CP_9964_elements(15) & timerDaemon_CP_9964_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3825_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/aggregated_phi_sample_ack
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(35) & timerDaemon_CP_9964_elements(17);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(32) & timerDaemon_CP_9964_elements(16);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(36) & timerDaemon_CP_9964_elements(18);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(9) & timerDaemon_CP_9964_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(9) & timerDaemon_CP_9964_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_9964_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	37 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_update_completed_
      -- 
    -- Element group timerDaemon_CP_9964_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_loopback_trigger
      -- 
    timerDaemon_CP_9964_elements(19) <= timerDaemon_CP_9964_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_loopback_sample_req_ps
      -- 
    phi_stmt_3820_loopback_sample_req_10003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3820_loopback_sample_req_10003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(20), ack => phi_stmt_3820_req_1); -- 
    -- Element group timerDaemon_CP_9964_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_entry_trigger
      -- 
    timerDaemon_CP_9964_elements(21) <= timerDaemon_CP_9964_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_entry_sample_req
      -- 
    phi_stmt_3820_entry_sample_req_10006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3820_entry_sample_req_10006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(22), ack => phi_stmt_3820_req_0); -- 
    -- Element group timerDaemon_CP_9964_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3820_phi_mux_ack_ps
      -- 
    phi_stmt_3820_phi_mux_ack_10009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3820_ack_0, ack => timerDaemon_CP_9964_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/type_cast_3823_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/type_cast_3823_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/type_cast_3823_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/type_cast_3823_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_9964_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/type_cast_3823_update_start_
      -- CP-element group 25: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/type_cast_3823_update_start__ps
      -- 
    -- Element group timerDaemon_CP_9964_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/type_cast_3823_update_completed__ps
      -- 
    timerDaemon_CP_9964_elements(26) <= timerDaemon_CP_9964_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/type_cast_3823_update_completed_
      -- 
    -- Element group timerDaemon_CP_9964_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_9964_elements(25), ack => timerDaemon_CP_9964_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_sample_start__ps
      -- 
    req_10030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(28), ack => nCOUNTER_3833_3824_buf_req_0); -- 
    -- Element group timerDaemon_CP_9964_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_Update/req
      -- CP-element group 29: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_update_start_
      -- CP-element group 29: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_update_start__ps
      -- 
    req_10035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(29), ack => nCOUNTER_3833_3824_buf_req_1); -- 
    -- Element group timerDaemon_CP_9964_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_sample_completed_
      -- 
    ack_10031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3833_3824_buf_ack_0, ack => timerDaemon_CP_9964_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/R_nCOUNTER_3824_Update/$exit
      -- 
    ack_10036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3833_3824_buf_ack_1, ack => timerDaemon_CP_9964_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3825_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(9) & timerDaemon_CP_9964_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_Sample/rr
      -- 
    rr_10049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_10049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(33), ack => RPIPE_timer_req_3827_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(11) & timerDaemon_CP_9964_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_update_start_
      -- CP-element group 34: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_Update/$entry
      -- 
    cr_10054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_10054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(34), ack => RPIPE_timer_req_3827_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(35) & timerDaemon_CP_9964_elements(13);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_Sample/ra
      -- 
    ra_10050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_3827_inst_ack_0, ack => timerDaemon_CP_9964_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/phi_stmt_3825_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/RPIPE_timer_req_3827_Update/$exit
      -- 
    ca_10055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_3827_inst_ack_1, ack => timerDaemon_CP_9964_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	18 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_sample_start_
      -- 
    req_10063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(37), ack => WPIPE_timer_resp_3835_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(36) & timerDaemon_CP_9964_elements(18) & timerDaemon_CP_9964_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_Update/req
      -- CP-element group 38: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_update_start_
      -- CP-element group 38: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_sample_completed_
      -- 
    ack_10064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_3835_inst_ack_0, ack => timerDaemon_CP_9964_elements(38)); -- 
    req_10068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_10068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9964_elements(38), ack => WPIPE_timer_resp_3835_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/WPIPE_timer_resp_3835_update_completed_
      -- 
    ack_10069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_3835_inst_ack_1, ack => timerDaemon_CP_9964_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_9964_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_9964_elements(9), ack => timerDaemon_CP_9964_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_3817/do_while_stmt_3818/do_while_stmt_3818_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9964_elements(39) & timerDaemon_CP_9964_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9964_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_3817/do_while_stmt_3818/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_3817/do_while_stmt_3818/loop_exit/ack
      -- 
    ack_10074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3818_branch_ack_0, ack => timerDaemon_CP_9964_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_3817/do_while_stmt_3818/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_3817/do_while_stmt_3818/loop_taken/ack
      -- 
    ack_10078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3818_branch_ack_1, ack => timerDaemon_CP_9964_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_3817/do_while_stmt_3818/$exit
      -- 
    timerDaemon_CP_9964_elements(44) <= timerDaemon_CP_9964_elements(3);
    timerDaemon_do_while_stmt_3818_terminator_10079: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_3818_terminator_10079", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_9964_elements(6),loop_continue => timerDaemon_CP_9964_elements(43),loop_terminate => timerDaemon_CP_9964_elements(42),loop_back => timerDaemon_CP_9964_elements(4),loop_exit => timerDaemon_CP_9964_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_3820_phi_seq_10037_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_9964_elements(21);
      timerDaemon_CP_9964_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_9964_elements(24);
      timerDaemon_CP_9964_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_9964_elements(26);
      timerDaemon_CP_9964_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_9964_elements(19);
      timerDaemon_CP_9964_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_9964_elements(30);
      timerDaemon_CP_9964_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_9964_elements(31);
      timerDaemon_CP_9964_elements(20) <= phi_mux_reqs(1);
      phi_stmt_3820_phi_seq_10037 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_3820_phi_seq_10037") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_9964_elements(11), 
          phi_sample_ack => timerDaemon_CP_9964_elements(17), 
          phi_update_req => timerDaemon_CP_9964_elements(13), 
          phi_update_ack => timerDaemon_CP_9964_elements(18), 
          phi_mux_ack => timerDaemon_CP_9964_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_9989_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_9964_elements(7);
        preds(1)  <= timerDaemon_CP_9964_elements(8);
        entry_tmerge_9989 : transition_merge -- 
          generic map(name => " entry_tmerge_9989")
          port map (preds => preds, symbol_out => timerDaemon_CP_9964_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_3820 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_3827_wire : std_logic_vector(0 downto 0);
    signal konst_3831_wire_constant : std_logic_vector(63 downto 0);
    signal konst_3839_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_3833 : std_logic_vector(63 downto 0);
    signal nCOUNTER_3833_3824_buffered : std_logic_vector(63 downto 0);
    signal req_3825 : std_logic_vector(0 downto 0);
    signal type_cast_3823_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_3831_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_3839_wire_constant <= "1";
    type_cast_3823_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_3820: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3823_wire_constant & nCOUNTER_3833_3824_buffered;
      req <= phi_stmt_3820_req_0 & phi_stmt_3820_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3820",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3820_ack_0,
          idata => idata,
          odata => COUNTER_3820,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3820
    nCOUNTER_3833_3824_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_3833_3824_buf_req_0;
      nCOUNTER_3833_3824_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_3833_3824_buf_req_1;
      nCOUNTER_3833_3824_buf_ack_1<= rack(0);
      nCOUNTER_3833_3824_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_3833_3824_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_3833,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_3833_3824_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_3825
    process(RPIPE_timer_req_3827_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_3827_wire(0 downto 0);
      req_3825 <= tmp_var; -- 
    end process;
    do_while_stmt_3818_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_3839_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3818_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3818_branch_req_0,
          ack0 => do_while_stmt_3818_branch_ack_0,
          ack1 => do_while_stmt_3818_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_3832_inst
    process(COUNTER_3820) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_3820, konst_3831_wire_constant, tmp_var);
      nCOUNTER_3833 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_3827_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_3827_inst_req_0;
      RPIPE_timer_req_3827_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_3827_inst_req_1;
      RPIPE_timer_req_3827_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_3827_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_3835_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_3835_inst_req_0;
      WPIPE_timer_resp_3835_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_3835_inst_req_1;
      WPIPE_timer_resp_3835_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_3825(0);
      data_in <= COUNTER_3820;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(27 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(127 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(27 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(127 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(20 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_row_in :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(47 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(47 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(47 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(63 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe4_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_num_chl :  std_logic_vector(15 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(79 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(79 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(63 downto 0);
  signal sendB_in_args    : std_logic_vector(63 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(63 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendModule
  component sendModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
      output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendModule
  signal sendModule_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendModule_tag_out   : std_logic_vector(1 downto 0);
  signal sendModule_start_req : std_logic;
  signal sendModule_start_ack : std_logic;
  signal sendModule_fin_req   : std_logic;
  signal sendModule_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe2
  signal input_pipe2_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe2
  signal input_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe3
  signal input_pipe3_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe3
  signal input_pipe3_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe4
  signal input_pipe4_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe4_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe4
  signal input_pipe4_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe4_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe2
  signal kernel_pipe2_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe2
  signal kernel_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe3
  signal kernel_pipe3_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe3
  signal kernel_pipe3_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe output_pipe
  signal output_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe output_pipe
  signal output_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_row_in <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 48,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      row_in => access_T_row_in,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(20 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 0),
      input_pipe2_pipe_write_req => input_pipe2_pipe_write_req(0 downto 0),
      input_pipe2_pipe_write_ack => input_pipe2_pipe_write_ack(0 downto 0),
      input_pipe2_pipe_write_data => input_pipe2_pipe_write_data(15 downto 0),
      input_pipe3_pipe_write_req => input_pipe3_pipe_write_req(0 downto 0),
      input_pipe3_pipe_write_ack => input_pipe3_pipe_write_ack(0 downto 0),
      input_pipe3_pipe_write_data => input_pipe3_pipe_write_data(15 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      input_pipe4_pipe_write_req => input_pipe4_pipe_write_req(0 downto 0),
      input_pipe4_pipe_write_ack => input_pipe4_pipe_write_ack(0 downto 0),
      input_pipe4_pipe_write_data => input_pipe4_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(27 downto 14),
      memory_space_0_sr_data => memory_space_0_sr_data(127 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(39 downto 20),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(20 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(7 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(1 downto 1),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(1 downto 1),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(31 downto 16),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(47 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(79 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(63 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe2_pipe_read_req => input_pipe2_pipe_read_req(0 downto 0),
      input_pipe2_pipe_read_ack => input_pipe2_pipe_read_ack(0 downto 0),
      input_pipe2_pipe_read_data => input_pipe2_pipe_read_data(15 downto 0),
      input_pipe3_pipe_read_req => input_pipe3_pipe_read_req(0 downto 0),
      input_pipe3_pipe_read_ack => input_pipe3_pipe_read_ack(0 downto 0),
      input_pipe3_pipe_read_data => input_pipe3_pipe_read_data(15 downto 0),
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      kernel_pipe2_pipe_read_req => kernel_pipe2_pipe_read_req(0 downto 0),
      kernel_pipe2_pipe_read_ack => kernel_pipe2_pipe_read_ack(0 downto 0),
      kernel_pipe2_pipe_read_data => kernel_pipe2_pipe_read_data(15 downto 0),
      kernel_pipe3_pipe_read_req => kernel_pipe3_pipe_read_req(0 downto 0),
      kernel_pipe3_pipe_read_ack => kernel_pipe3_pipe_read_ack(0 downto 0),
      kernel_pipe3_pipe_read_data => kernel_pipe3_pipe_read_data(15 downto 0),
      input_pipe4_pipe_read_req => input_pipe4_pipe_read_req(0 downto 0),
      input_pipe4_pipe_read_ack => input_pipe4_pipe_read_ack(0 downto 0),
      input_pipe4_pipe_read_data => input_pipe4_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(1 downto 1),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(1 downto 1),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(15 downto 8),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(0 downto 0),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(0 downto 0),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(79 downto 16);
  loadKernelChannel_num_chl <= loadKernelChannel_in_args(15 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 80,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      num_chl => loadKernelChannel_num_chl,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(1 downto 1),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(1 downto 1),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(15 downto 8),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(0 downto 0),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(0 downto 0),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(15 downto 0),
      kernel_pipe3_pipe_write_req => kernel_pipe3_pipe_write_req(0 downto 0),
      kernel_pipe3_pipe_write_ack => kernel_pipe3_pipe_write_ack(0 downto 0),
      kernel_pipe3_pipe_write_data => kernel_pipe3_pipe_write_data(15 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(15 downto 0),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(63 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module sendModule
  sendModule_instance:sendModule-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendModule_start_req,
      start_ack => sendModule_start_ack,
      fin_req => sendModule_fin_req,
      fin_ack => sendModule_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      output_pipe_pipe_read_req => output_pipe_pipe_read_req(1 downto 0),
      output_pipe_pipe_read_ack => output_pipe_pipe_read_ack(1 downto 0),
      output_pipe_pipe_read_data => output_pipe_pipe_read_data(31 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(7 downto 0),
      tag_in => sendModule_tag_in,
      tag_out => sendModule_tag_out-- 
    ); -- 
  -- module will be run forever 
  sendModule_tag_in <= (others => '0');
  sendModule_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => sendModule_start_req, start_ack => sendModule_start_ack,  fin_req => sendModule_fin_req,  fin_ack => sendModule_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe2_pipe_read_req,
      read_ack => input_pipe2_pipe_read_ack,
      read_data => input_pipe2_pipe_read_data,
      write_req => input_pipe2_pipe_write_req,
      write_ack => input_pipe2_pipe_write_ack,
      write_data => input_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe3_pipe_read_req,
      read_ack => input_pipe3_pipe_read_ack,
      read_data => input_pipe3_pipe_read_data,
      write_req => input_pipe3_pipe_write_req,
      write_ack => input_pipe3_pipe_write_ack,
      write_data => input_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe4",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe4_pipe_read_req,
      read_ack => input_pipe4_pipe_read_ack,
      read_data => input_pipe4_pipe_read_data,
      write_req => input_pipe4_pipe_write_req,
      write_ack => input_pipe4_pipe_write_ack,
      write_data => input_pipe4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe2_pipe_read_req,
      read_ack => kernel_pipe2_pipe_read_ack,
      read_data => kernel_pipe2_pipe_read_data,
      write_req => kernel_pipe2_pipe_write_req,
      write_ack => kernel_pipe2_pipe_write_ack,
      write_data => kernel_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe3_pipe_read_req,
      read_ack => kernel_pipe3_pipe_read_ack,
      read_data => kernel_pipe3_pipe_read_data,
      write_req => kernel_pipe3_pipe_write_req,
      write_ack => kernel_pipe3_pipe_write_ack,
      write_data => kernel_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe output_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 10 --
    )
    port map( -- 
      read_req => output_pipe_pipe_read_req,
      read_ack => output_pipe_pipe_read_ack,
      read_data => output_pipe_pipe_read_data,
      write_req => output_pipe_pipe_write_req,
      write_ack => output_pipe_pipe_write_ack,
      write_data => output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 11 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 2,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 4,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
