-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant Kernel_base_address : std_logic_vector(18 downto 0) := "0000000000000000000";
  constant Tensor0_base_address : std_logic_vector(18 downto 0) := "0000000000000000000";
  constant Tensor1_base_address : std_logic_vector(19 downto 0) := "00000000000000000000";
  constant Tensor2_base_address : std_logic_vector(18 downto 0) := "0000000000000000000";
  constant Tensor3_base_address : std_logic_vector(17 downto 0) := "000000000000000000";
  constant Tensor4_base_address : std_logic_vector(16 downto 0) := "00000000000000000";
  -- 
end package ahir_system_global_package;
