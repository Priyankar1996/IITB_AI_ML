-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_3606_start: Boolean;
  signal convTranspose_CP_3606_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1225_call_req_0 : boolean;
  signal call_stmt_1225_call_ack_0 : boolean;
  signal call_stmt_1225_call_req_1 : boolean;
  signal call_stmt_1225_call_ack_1 : boolean;
  signal WPIPE_Block0_start_1227_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1227_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1227_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1227_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1230_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1230_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1230_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1230_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1233_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1233_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1233_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1233_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1236_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1236_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1236_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1236_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1241_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1241_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1241_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1241_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1244_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1244_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1244_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1244_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1247_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1247_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1247_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1247_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1250_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1250_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1250_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1250_inst_ack_1 : boolean;
  signal call_stmt_1253_call_req_0 : boolean;
  signal call_stmt_1253_call_ack_0 : boolean;
  signal call_stmt_1253_call_req_1 : boolean;
  signal call_stmt_1253_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_3606_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3606_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_3606_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3606_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_3606: Block -- control-path 
    signal convTranspose_CP_3606_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    convTranspose_CP_3606_elements(0) <= convTranspose_CP_3606_start;
    convTranspose_CP_3606_symbol <= convTranspose_CP_3606_elements(22);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1223/$entry
      -- CP-element group 0: 	 branch_block_stmt_1223/branch_block_stmt_1223__entry__
      -- CP-element group 0: 	 branch_block_stmt_1223/call_stmt_1225__entry__
      -- CP-element group 0: 	 branch_block_stmt_1223/call_stmt_1225/$entry
      -- CP-element group 0: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_Update/ccr
      -- 
    crr_3634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(0), ack => call_stmt_1225_call_req_0); -- 
    ccr_3639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(0), ack => call_stmt_1225_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_Sample/cra
      -- 
    cra_3635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1225_call_ack_0, ack => convTranspose_CP_3606_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (19) 
      -- CP-element group 2: 	 branch_block_stmt_1223/call_stmt_1225__exit__
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238__entry__
      -- CP-element group 2: 	 branch_block_stmt_1223/call_stmt_1225/$exit
      -- CP-element group 2: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1223/call_stmt_1225/call_stmt_1225_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/$entry
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_Sample/req
      -- 
    cca_3640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1225_call_ack_1, ack => convTranspose_CP_3606_elements(2)); -- 
    req_3651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(2), ack => WPIPE_Block0_start_1227_inst_req_0); -- 
    req_3665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(2), ack => WPIPE_Block1_start_1230_inst_req_0); -- 
    req_3679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(2), ack => WPIPE_Block2_start_1233_inst_req_0); -- 
    req_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(2), ack => WPIPE_Block3_start_1236_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_Update/req
      -- 
    ack_3652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1227_inst_ack_0, ack => convTranspose_CP_3606_elements(3)); -- 
    req_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(3), ack => WPIPE_Block0_start_1227_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	11 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block0_start_1227_Update/ack
      -- 
    ack_3657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1227_inst_ack_1, ack => convTranspose_CP_3606_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_Update/req
      -- 
    ack_3666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1230_inst_ack_0, ack => convTranspose_CP_3606_elements(5)); -- 
    req_3670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(5), ack => WPIPE_Block1_start_1230_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	11 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block1_start_1230_Update/ack
      -- 
    ack_3671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1230_inst_ack_1, ack => convTranspose_CP_3606_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_Update/req
      -- 
    ack_3680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1233_inst_ack_0, ack => convTranspose_CP_3606_elements(7)); -- 
    req_3684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(7), ack => WPIPE_Block2_start_1233_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block2_start_1233_Update/ack
      -- 
    ack_3685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1233_inst_ack_1, ack => convTranspose_CP_3606_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_Update/req
      -- 
    ack_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1236_inst_ack_0, ack => convTranspose_CP_3606_elements(9)); -- 
    req_3698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(9), ack => WPIPE_Block3_start_1236_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/WPIPE_Block3_start_1236_Update/ack
      -- 
    ack_3699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1236_inst_ack_1, ack => convTranspose_CP_3606_elements(10)); -- 
    -- CP-element group 11:  join  fork  transition  place  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	10 
    -- CP-element group 11: 	4 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	18 
    -- CP-element group 11:  members (16) 
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238__exit__
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251__entry__
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1229_to_assign_stmt_1238/$exit
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/$entry
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_Sample/rr
      -- 
    rr_3710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(11), ack => RPIPE_Block0_done_1241_inst_req_0); -- 
    rr_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(11), ack => RPIPE_Block1_done_1244_inst_req_0); -- 
    rr_3738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(11), ack => RPIPE_Block2_done_1247_inst_req_0); -- 
    rr_3752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(11), ack => RPIPE_Block3_done_1250_inst_req_0); -- 
    convTranspose_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_3606_elements(8) & convTranspose_CP_3606_elements(6) & convTranspose_CP_3606_elements(10) & convTranspose_CP_3606_elements(4);
      gj_convTranspose_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3606_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_Update/cr
      -- 
    ra_3711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1241_inst_ack_0, ack => convTranspose_CP_3606_elements(12)); -- 
    cr_3715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(12), ack => RPIPE_Block0_done_1241_inst_req_1); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	20 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block0_done_1241_Update/ca
      -- 
    ca_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1241_inst_ack_1, ack => convTranspose_CP_3606_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_Update/cr
      -- 
    ra_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1244_inst_ack_0, ack => convTranspose_CP_3606_elements(14)); -- 
    cr_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(14), ack => RPIPE_Block1_done_1244_inst_req_1); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block1_done_1244_Update/ca
      -- 
    ca_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1244_inst_ack_1, ack => convTranspose_CP_3606_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_Update/cr
      -- 
    ra_3739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1247_inst_ack_0, ack => convTranspose_CP_3606_elements(16)); -- 
    cr_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(16), ack => RPIPE_Block2_done_1247_inst_req_1); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	20 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block2_done_1247_Update/ca
      -- 
    ca_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1247_inst_ack_1, ack => convTranspose_CP_3606_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_Update/cr
      -- 
    ra_3753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1250_inst_ack_0, ack => convTranspose_CP_3606_elements(18)); -- 
    cr_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(18), ack => RPIPE_Block3_done_1250_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/RPIPE_Block3_done_1250_Update/ca
      -- 
    ca_3758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1250_inst_ack_1, ack => convTranspose_CP_3606_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  place  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	19 
    -- CP-element group 20: 	13 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (10) 
      -- CP-element group 20: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251__exit__
      -- CP-element group 20: 	 branch_block_stmt_1223/call_stmt_1253__entry__
      -- CP-element group 20: 	 branch_block_stmt_1223/assign_stmt_1242_to_assign_stmt_1251/$exit
      -- CP-element group 20: 	 branch_block_stmt_1223/call_stmt_1253/$entry
      -- CP-element group 20: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_Sample/crr
      -- CP-element group 20: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_Update/ccr
      -- 
    crr_3769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(20), ack => call_stmt_1253_call_req_0); -- 
    ccr_3774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3606_elements(20), ack => call_stmt_1253_call_req_1); -- 
    convTranspose_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTranspose_CP_3606_elements(15) & convTranspose_CP_3606_elements(17) & convTranspose_CP_3606_elements(19) & convTranspose_CP_3606_elements(13);
      gj_convTranspose_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3606_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_Sample/cra
      -- 
    cra_3770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1253_call_ack_0, ack => convTranspose_CP_3606_elements(21)); -- 
    -- CP-element group 22:  transition  place  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (16) 
      -- CP-element group 22: 	 $exit
      -- CP-element group 22: 	 branch_block_stmt_1223/$exit
      -- CP-element group 22: 	 branch_block_stmt_1223/branch_block_stmt_1223__exit__
      -- CP-element group 22: 	 branch_block_stmt_1223/call_stmt_1253__exit__
      -- CP-element group 22: 	 branch_block_stmt_1223/return__
      -- CP-element group 22: 	 branch_block_stmt_1223/merge_stmt_1255__exit__
      -- CP-element group 22: 	 branch_block_stmt_1223/call_stmt_1253/$exit
      -- CP-element group 22: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1223/call_stmt_1253/call_stmt_1253_Update/cca
      -- CP-element group 22: 	 branch_block_stmt_1223/return___PhiReq/$entry
      -- CP-element group 22: 	 branch_block_stmt_1223/return___PhiReq/$exit
      -- CP-element group 22: 	 branch_block_stmt_1223/merge_stmt_1255_PhiReqMerge
      -- CP-element group 22: 	 branch_block_stmt_1223/merge_stmt_1255_PhiAck/$entry
      -- CP-element group 22: 	 branch_block_stmt_1223/merge_stmt_1255_PhiAck/$exit
      -- CP-element group 22: 	 branch_block_stmt_1223/merge_stmt_1255_PhiAck/dummy
      -- 
    cca_3775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1253_call_ack_1, ack => convTranspose_CP_3606_elements(22)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call11_1251 : std_logic_vector(15 downto 0);
    signal call5_1242 : std_logic_vector(15 downto 0);
    signal call7_1245 : std_logic_vector(15 downto 0);
    signal call9_1248 : std_logic_vector(15 downto 0);
    signal call_1225 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    -- shared inport operator group (0) : RPIPE_Block0_done_1241_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1241_inst_req_0;
      RPIPE_Block0_done_1241_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1241_inst_req_1;
      RPIPE_Block0_done_1241_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call5_1242 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1244_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1244_inst_req_0;
      RPIPE_Block1_done_1244_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1244_inst_req_1;
      RPIPE_Block1_done_1244_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call7_1245 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1247_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1247_inst_req_0;
      RPIPE_Block2_done_1247_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1247_inst_req_1;
      RPIPE_Block2_done_1247_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call9_1248 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1250_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1250_inst_req_0;
      RPIPE_Block3_done_1250_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1250_inst_req_1;
      RPIPE_Block3_done_1250_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call11_1251 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_start_1227_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_start_1227_inst_req_0;
      WPIPE_Block0_start_1227_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_start_1227_inst_req_1;
      WPIPE_Block0_start_1227_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1225;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1230_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_start_1230_inst_req_0;
      WPIPE_Block1_start_1230_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_start_1230_inst_req_1;
      WPIPE_Block1_start_1230_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1225;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1233_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_start_1233_inst_req_0;
      WPIPE_Block2_start_1233_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_start_1233_inst_req_1;
      WPIPE_Block2_start_1233_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1225;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1236_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_start_1236_inst_req_0;
      WPIPE_Block3_start_1236_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_start_1236_inst_req_1;
      WPIPE_Block3_start_1236_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1225;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1225_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1225_call_req_0;
      call_stmt_1225_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1225_call_req_1;
      call_stmt_1225_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1225 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1253_call 
    sendOutput_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1253_call_req_0;
      call_stmt_1253_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1253_call_req_1;
      call_stmt_1253_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3784_start: Boolean;
  signal convTransposeA_CP_3784_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1321_load_0_ack_1 : boolean;
  signal LOAD_padding_1311_load_0_ack_0 : boolean;
  signal ptr_deref_1286_load_0_ack_1 : boolean;
  signal LOAD_padding_1311_load_0_ack_1 : boolean;
  signal ptr_deref_1321_load_0_req_1 : boolean;
  signal LOAD_padding_1311_load_0_req_0 : boolean;
  signal ptr_deref_1274_load_0_req_1 : boolean;
  signal ptr_deref_1274_load_0_ack_1 : boolean;
  signal RPIPE_Block0_start_1261_inst_ack_0 : boolean;
  signal ptr_deref_1308_load_0_req_0 : boolean;
  signal ptr_deref_1308_load_0_ack_0 : boolean;
  signal ptr_deref_1286_load_0_req_1 : boolean;
  signal RPIPE_Block0_start_1261_inst_req_0 : boolean;
  signal ptr_deref_1296_load_0_req_0 : boolean;
  signal ptr_deref_1296_load_0_ack_0 : boolean;
  signal LOAD_padding_1311_load_0_req_1 : boolean;
  signal ptr_deref_1296_load_0_req_1 : boolean;
  signal RPIPE_Block0_start_1261_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1261_inst_ack_1 : boolean;
  signal ptr_deref_1296_load_0_ack_1 : boolean;
  signal ptr_deref_1286_load_0_req_0 : boolean;
  signal ptr_deref_1286_load_0_ack_0 : boolean;
  signal ptr_deref_1308_load_0_req_1 : boolean;
  signal ptr_deref_1321_load_0_ack_0 : boolean;
  signal ptr_deref_1308_load_0_ack_1 : boolean;
  signal ptr_deref_1333_load_0_req_0 : boolean;
  signal ptr_deref_1333_load_0_ack_0 : boolean;
  signal ptr_deref_1321_load_0_req_0 : boolean;
  signal ptr_deref_1274_load_0_ack_0 : boolean;
  signal ptr_deref_1274_load_0_req_0 : boolean;
  signal ptr_deref_1333_load_0_req_1 : boolean;
  signal ptr_deref_1333_load_0_ack_1 : boolean;
  signal ptr_deref_1345_load_0_req_0 : boolean;
  signal ptr_deref_1345_load_0_ack_0 : boolean;
  signal ptr_deref_1345_load_0_req_1 : boolean;
  signal ptr_deref_1345_load_0_ack_1 : boolean;
  signal ptr_deref_1357_load_0_req_0 : boolean;
  signal ptr_deref_1357_load_0_ack_0 : boolean;
  signal ptr_deref_1357_load_0_req_1 : boolean;
  signal ptr_deref_1357_load_0_ack_1 : boolean;
  signal type_cast_1361_inst_req_0 : boolean;
  signal type_cast_1361_inst_ack_0 : boolean;
  signal type_cast_1361_inst_req_1 : boolean;
  signal type_cast_1361_inst_ack_1 : boolean;
  signal type_cast_1365_inst_req_0 : boolean;
  signal type_cast_1365_inst_ack_0 : boolean;
  signal type_cast_1365_inst_req_1 : boolean;
  signal type_cast_1365_inst_ack_1 : boolean;
  signal ptr_deref_1383_load_0_req_0 : boolean;
  signal ptr_deref_1383_load_0_ack_0 : boolean;
  signal ptr_deref_1383_load_0_req_1 : boolean;
  signal ptr_deref_1383_load_0_ack_1 : boolean;
  signal type_cast_1387_inst_req_0 : boolean;
  signal type_cast_1387_inst_ack_0 : boolean;
  signal type_cast_1387_inst_req_1 : boolean;
  signal type_cast_1387_inst_ack_1 : boolean;
  signal type_cast_1512_inst_req_0 : boolean;
  signal type_cast_1512_inst_ack_0 : boolean;
  signal type_cast_1512_inst_req_1 : boolean;
  signal type_cast_1512_inst_ack_1 : boolean;
  signal array_obj_ref_1524_index_offset_req_0 : boolean;
  signal array_obj_ref_1524_index_offset_ack_0 : boolean;
  signal array_obj_ref_1524_index_offset_req_1 : boolean;
  signal array_obj_ref_1524_index_offset_ack_1 : boolean;
  signal addr_of_1525_final_reg_req_0 : boolean;
  signal addr_of_1525_final_reg_ack_0 : boolean;
  signal addr_of_1525_final_reg_req_1 : boolean;
  signal addr_of_1525_final_reg_ack_1 : boolean;
  signal ptr_deref_1529_load_0_req_0 : boolean;
  signal ptr_deref_1529_load_0_ack_0 : boolean;
  signal ptr_deref_1529_load_0_req_1 : boolean;
  signal ptr_deref_1529_load_0_ack_1 : boolean;
  signal type_cast_1533_inst_req_0 : boolean;
  signal type_cast_1533_inst_ack_0 : boolean;
  signal type_cast_1533_inst_req_1 : boolean;
  signal type_cast_1533_inst_ack_1 : boolean;
  signal array_obj_ref_1545_index_offset_req_0 : boolean;
  signal array_obj_ref_1545_index_offset_ack_0 : boolean;
  signal array_obj_ref_1545_index_offset_req_1 : boolean;
  signal array_obj_ref_1545_index_offset_ack_1 : boolean;
  signal addr_of_1546_final_reg_req_0 : boolean;
  signal addr_of_1546_final_reg_ack_0 : boolean;
  signal addr_of_1546_final_reg_req_1 : boolean;
  signal addr_of_1546_final_reg_ack_1 : boolean;
  signal ptr_deref_1549_store_0_req_0 : boolean;
  signal ptr_deref_1549_store_0_ack_0 : boolean;
  signal ptr_deref_1549_store_0_req_1 : boolean;
  signal ptr_deref_1549_store_0_ack_1 : boolean;
  signal type_cast_1554_inst_req_0 : boolean;
  signal type_cast_1554_inst_ack_0 : boolean;
  signal type_cast_1554_inst_req_1 : boolean;
  signal type_cast_1554_inst_ack_1 : boolean;
  signal if_stmt_1567_branch_req_0 : boolean;
  signal if_stmt_1567_branch_ack_1 : boolean;
  signal if_stmt_1567_branch_ack_0 : boolean;
  signal type_cast_1590_inst_req_0 : boolean;
  signal type_cast_1590_inst_ack_0 : boolean;
  signal type_cast_1590_inst_req_1 : boolean;
  signal type_cast_1590_inst_ack_1 : boolean;
  signal type_cast_1599_inst_req_0 : boolean;
  signal type_cast_1599_inst_ack_0 : boolean;
  signal type_cast_1599_inst_req_1 : boolean;
  signal type_cast_1599_inst_ack_1 : boolean;
  signal type_cast_1615_inst_req_0 : boolean;
  signal type_cast_1615_inst_ack_0 : boolean;
  signal type_cast_1615_inst_req_1 : boolean;
  signal type_cast_1615_inst_ack_1 : boolean;
  signal if_stmt_1622_branch_req_0 : boolean;
  signal if_stmt_1622_branch_ack_1 : boolean;
  signal if_stmt_1622_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1630_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1630_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1630_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1630_inst_ack_1 : boolean;
  signal phi_stmt_1419_req_0 : boolean;
  signal phi_stmt_1426_req_0 : boolean;
  signal type_cast_1425_inst_req_0 : boolean;
  signal type_cast_1425_inst_ack_0 : boolean;
  signal type_cast_1425_inst_req_1 : boolean;
  signal type_cast_1425_inst_ack_1 : boolean;
  signal phi_stmt_1419_req_1 : boolean;
  signal type_cast_1432_inst_req_0 : boolean;
  signal type_cast_1432_inst_ack_0 : boolean;
  signal type_cast_1432_inst_req_1 : boolean;
  signal type_cast_1432_inst_ack_1 : boolean;
  signal phi_stmt_1426_req_1 : boolean;
  signal phi_stmt_1419_ack_0 : boolean;
  signal phi_stmt_1426_ack_0 : boolean;
  signal type_cast_1492_inst_req_0 : boolean;
  signal type_cast_1492_inst_ack_0 : boolean;
  signal type_cast_1492_inst_req_1 : boolean;
  signal type_cast_1492_inst_ack_1 : boolean;
  signal phi_stmt_1486_req_1 : boolean;
  signal phi_stmt_1486_req_0 : boolean;
  signal phi_stmt_1486_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3784_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3784_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3784_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3784_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3784: Block -- control-path 
    signal convTransposeA_CP_3784_elements: BooleanArray(81 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3784_elements(0) <= convTransposeA_CP_3784_start;
    convTransposeA_CP_3784_symbol <= convTransposeA_CP_3784_elements(61);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1259/assign_stmt_1262__entry__
      -- CP-element group 0: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1259/assign_stmt_1262/$entry
      -- CP-element group 0: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1259/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1259/branch_block_stmt_1259__entry__
      -- 
    rr_3832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(0), ack => RPIPE_Block0_start_1261_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_sample_completed_
      -- 
    ra_3833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1261_inst_ack_0, ack => convTransposeA_CP_3784_elements(1)); -- 
    cr_3837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(1), ack => RPIPE_Block0_start_1261_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1262__exit__
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416__entry__
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1262/RPIPE_Block0_start_1261_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1262/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_Update/cr
      -- 
    ca_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1261_inst_ack_1, ack => convTransposeA_CP_3784_elements(2)); -- 
    cr_4118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1321_load_0_req_1); -- 
    rr_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => LOAD_padding_1311_load_0_req_0); -- 
    cr_3885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1274_load_0_req_1); -- 
    rr_4024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1308_load_0_req_0); -- 
    cr_3935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1286_load_0_req_1); -- 
    rr_3974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1296_load_0_req_0); -- 
    cr_4068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => LOAD_padding_1311_load_0_req_1); -- 
    cr_3985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1296_load_0_req_1); -- 
    rr_3924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1286_load_0_req_0); -- 
    cr_4035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1308_load_0_req_1); -- 
    rr_4157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1333_load_0_req_0); -- 
    rr_4107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1321_load_0_req_0); -- 
    rr_3874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1274_load_0_req_0); -- 
    cr_4168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1333_load_0_req_1); -- 
    rr_4207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1345_load_0_req_0); -- 
    cr_4218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1345_load_0_req_1); -- 
    rr_4257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1357_load_0_req_0); -- 
    cr_4268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1357_load_0_req_1); -- 
    cr_4287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => type_cast_1361_inst_req_1); -- 
    cr_4301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => type_cast_1365_inst_req_1); -- 
    rr_4335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1383_load_0_req_0); -- 
    cr_4346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => ptr_deref_1383_load_0_req_1); -- 
    cr_4365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(2), ack => type_cast_1387_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Sample/word_access_start/word_0/ra
      -- 
    ra_3875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1274_load_0_ack_0, ack => convTransposeA_CP_3784_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	21 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/ptr_deref_1274_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/ptr_deref_1274_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/ptr_deref_1274_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/ptr_deref_1274_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1274_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_Sample/rr
      -- 
    ca_3886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1274_load_0_ack_1, ack => convTransposeA_CP_3784_elements(4)); -- 
    rr_4282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(4), ack => type_cast_1361_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Sample/word_access_start/word_0/ra
      -- 
    ra_3925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1286_load_0_ack_0, ack => convTransposeA_CP_3784_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/ptr_deref_1286_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/ptr_deref_1286_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/ptr_deref_1286_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/ptr_deref_1286_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1286_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_Sample/rr
      -- 
    ca_3936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1286_load_0_ack_1, ack => convTransposeA_CP_3784_elements(6)); -- 
    rr_4296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(6), ack => type_cast_1365_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_sample_completed_
      -- 
    ra_3975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1296_load_0_ack_0, ack => convTransposeA_CP_3784_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	29 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/ptr_deref_1296_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/ptr_deref_1296_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/ptr_deref_1296_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1296_Update/ptr_deref_1296_Merge/merge_ack
      -- 
    ca_3986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1296_load_0_ack_1, ack => convTransposeA_CP_3784_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_sample_completed_
      -- 
    ra_4025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1308_load_0_ack_0, ack => convTransposeA_CP_3784_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/ptr_deref_1308_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/ptr_deref_1308_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/ptr_deref_1308_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/ptr_deref_1308_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1308_Update/word_access_complete/word_0/ca
      -- 
    ca_4036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1308_load_0_ack_1, ack => convTransposeA_CP_3784_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Sample/word_access_start/word_0/ra
      -- CP-element group 11: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Sample/word_access_start/word_0/$exit
      -- 
    ra_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1311_load_0_ack_0, ack => convTransposeA_CP_3784_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/LOAD_padding_1311_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/LOAD_padding_1311_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/LOAD_padding_1311_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/LOAD_padding_1311_Update/LOAD_padding_1311_Merge/merge_req
      -- 
    ca_4069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1311_load_0_ack_1, ack => convTransposeA_CP_3784_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Sample/word_access_start/word_0/$exit
      -- 
    ra_4108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1321_load_0_ack_0, ack => convTransposeA_CP_3784_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	29 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/ptr_deref_1321_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/ptr_deref_1321_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/ptr_deref_1321_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/ptr_deref_1321_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1321_update_completed_
      -- 
    ca_4119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1321_load_0_ack_1, ack => convTransposeA_CP_3784_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Sample/word_access_start/word_0/ra
      -- 
    ra_4158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1333_load_0_ack_0, ack => convTransposeA_CP_3784_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/ptr_deref_1333_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/ptr_deref_1333_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/ptr_deref_1333_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1333_Update/ptr_deref_1333_Merge/merge_ack
      -- 
    ca_4169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1333_load_0_ack_1, ack => convTransposeA_CP_3784_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Sample/word_access_start/word_0/ra
      -- 
    ra_4208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1345_load_0_ack_0, ack => convTransposeA_CP_3784_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	29 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/ptr_deref_1345_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/ptr_deref_1345_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/ptr_deref_1345_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1345_Update/ptr_deref_1345_Merge/merge_ack
      -- 
    ca_4219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1345_load_0_ack_1, ack => convTransposeA_CP_3784_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Sample/word_access_start/word_0/ra
      -- 
    ra_4258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_load_0_ack_0, ack => convTransposeA_CP_3784_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/ptr_deref_1357_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/ptr_deref_1357_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/ptr_deref_1357_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1357_Update/ptr_deref_1357_Merge/merge_ack
      -- 
    ca_4269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1357_load_0_ack_1, ack => convTransposeA_CP_3784_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	4 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_Sample/ra
      -- 
    ra_4283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_0, ack => convTransposeA_CP_3784_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1361_Update/ca
      -- 
    ca_4288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_1, ack => convTransposeA_CP_3784_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	6 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_Sample/ra
      -- 
    ra_4297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1365_inst_ack_0, ack => convTransposeA_CP_3784_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1365_Update/ca
      -- 
    ca_4302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1365_inst_ack_1, ack => convTransposeA_CP_3784_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Sample/word_access_start/word_0/ra
      -- 
    ra_4336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1383_load_0_ack_0, ack => convTransposeA_CP_3784_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (12) 
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/ptr_deref_1383_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/ptr_deref_1383_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/ptr_deref_1383_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/ptr_deref_1383_Update/ptr_deref_1383_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_Sample/rr
      -- 
    ca_4347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1383_load_0_ack_1, ack => convTransposeA_CP_3784_elements(26)); -- 
    rr_4360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(26), ack => type_cast_1387_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_Sample/ra
      -- 
    ra_4361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1387_inst_ack_0, ack => convTransposeA_CP_3784_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/type_cast_1387_Update/ca
      -- 
    ca_4366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1387_inst_ack_1, ack => convTransposeA_CP_3784_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	14 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	18 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	8 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	62 
    -- CP-element group 29: 	63 
    -- CP-element group 29:  members (8) 
      -- CP-element group 29: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416__exit__
      -- CP-element group 29: 	 branch_block_stmt_1259/assign_stmt_1271_to_assign_stmt_1416/$exit
      -- CP-element group 29: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/$entry
      -- CP-element group 29: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/$entry
      -- CP-element group 29: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/$entry
      -- 
    convTransposeA_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(20) & convTransposeA_CP_3784_elements(22) & convTransposeA_CP_3784_elements(24) & convTransposeA_CP_3784_elements(10) & convTransposeA_CP_3784_elements(12) & convTransposeA_CP_3784_elements(14) & convTransposeA_CP_3784_elements(16) & convTransposeA_CP_3784_elements(18) & convTransposeA_CP_3784_elements(28) & convTransposeA_CP_3784_elements(8);
      gj_convTransposeA_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	81 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_Sample/ra
      -- 
    ra_4381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1512_inst_ack_0, ack => convTransposeA_CP_3784_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	81 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (16) 
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_resized_1
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_scaled_1
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_computed_1
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_resize_1/$entry
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_resize_1/$exit
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_resize_1/index_resize_req
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_resize_1/index_resize_ack
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_scale_1/$entry
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_scale_1/$exit
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_scale_1/scale_rename_req
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_index_scale_1/scale_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_Sample/req
      -- 
    ca_4386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1512_inst_ack_1, ack => convTransposeA_CP_3784_elements(31)); -- 
    req_4411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(31), ack => array_obj_ref_1524_index_offset_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	49 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_sample_complete
      -- CP-element group 32: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_Sample/ack
      -- 
    ack_4412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1524_index_offset_ack_0, ack => convTransposeA_CP_3784_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	81 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (11) 
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_root_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_offset_calculated
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_Update/ack
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_base_plus_offset/$entry
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_base_plus_offset/$exit
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_base_plus_offset/sum_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_request/$entry
      -- CP-element group 33: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_request/req
      -- 
    ack_4417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1524_index_offset_ack_1, ack => convTransposeA_CP_3784_elements(33)); -- 
    req_4426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(33), ack => addr_of_1525_final_reg_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_request/$exit
      -- CP-element group 34: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_request/ack
      -- 
    ack_4427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1525_final_reg_ack_0, ack => convTransposeA_CP_3784_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	81 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (24) 
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_complete/ack
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_word_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_address_resized
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_addr_resize/$entry
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_addr_resize/$exit
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_word_addrgen/$entry
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_word_addrgen/$exit
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_word_addrgen/root_register_req
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_word_addrgen/root_register_ack
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Sample/word_access_start/$entry
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Sample/word_access_start/word_0/$entry
      -- CP-element group 35: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Sample/word_access_start/word_0/rr
      -- 
    ack_4432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1525_final_reg_ack_1, ack => convTransposeA_CP_3784_elements(35)); -- 
    rr_4465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(35), ack => ptr_deref_1529_load_0_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Sample/word_access_start/$exit
      -- CP-element group 36: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Sample/word_access_start/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Sample/word_access_start/word_0/ra
      -- 
    ra_4466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_load_0_ack_0, ack => convTransposeA_CP_3784_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	81 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	44 
    -- CP-element group 37:  members (9) 
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/word_access_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/word_access_complete/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/word_access_complete/word_0/ca
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/ptr_deref_1529_Merge/$entry
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/ptr_deref_1529_Merge/$exit
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/ptr_deref_1529_Merge/merge_req
      -- CP-element group 37: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/ptr_deref_1529_Merge/merge_ack
      -- 
    ca_4477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1529_load_0_ack_1, ack => convTransposeA_CP_3784_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	81 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_Sample/ra
      -- 
    ra_4491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1533_inst_ack_0, ack => convTransposeA_CP_3784_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	81 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (16) 
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_resized_1
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_scaled_1
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_computed_1
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_resize_1/$entry
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_resize_1/$exit
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_resize_1/index_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_resize_1/index_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_scale_1/$entry
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_scale_1/$exit
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_scale_1/scale_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_index_scale_1/scale_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_Sample/req
      -- 
    ca_4496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1533_inst_ack_1, ack => convTransposeA_CP_3784_elements(39)); -- 
    req_4521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(39), ack => array_obj_ref_1545_index_offset_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_sample_complete
      -- CP-element group 40: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_Sample/ack
      -- 
    ack_4522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1545_index_offset_ack_0, ack => convTransposeA_CP_3784_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	81 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (11) 
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_offset_calculated
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_request/$entry
      -- CP-element group 41: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_request/req
      -- 
    ack_4527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1545_index_offset_ack_1, ack => convTransposeA_CP_3784_elements(41)); -- 
    req_4536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(41), ack => addr_of_1546_final_reg_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_request/$exit
      -- CP-element group 42: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_request/ack
      -- 
    ack_4537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1546_final_reg_ack_0, ack => convTransposeA_CP_3784_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	81 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (19) 
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_complete/ack
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_word_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_address_resized
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_addr_resize/$entry
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_addr_resize/$exit
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_addr_resize/base_resize_req
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_addr_resize/base_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_word_addrgen/$entry
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_word_addrgen/$exit
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_word_addrgen/root_register_req
      -- CP-element group 43: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_word_addrgen/root_register_ack
      -- 
    ack_4542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1546_final_reg_ack_1, ack => convTransposeA_CP_3784_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	37 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/ptr_deref_1549_Split/$entry
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/ptr_deref_1549_Split/$exit
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/ptr_deref_1549_Split/split_req
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/ptr_deref_1549_Split/split_ack
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/word_access_start/word_0/rr
      -- 
    rr_4580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(44), ack => ptr_deref_1549_store_0_req_0); -- 
    convTransposeA_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(37) & convTransposeA_CP_3784_elements(43);
      gj_convTransposeA_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Sample/word_access_start/word_0/ra
      -- 
    ra_4581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1549_store_0_ack_0, ack => convTransposeA_CP_3784_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	81 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Update/word_access_complete/word_0/ca
      -- 
    ca_4592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1549_store_0_ack_1, ack => convTransposeA_CP_3784_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	81 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_Sample/ra
      -- 
    ra_4601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1554_inst_ack_0, ack => convTransposeA_CP_3784_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	81 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_Update/ca
      -- 
    ca_4606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1554_inst_ack_1, ack => convTransposeA_CP_3784_elements(48)); -- 
    -- CP-element group 49:  branch  join  transition  place  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	32 
    -- CP-element group 49: 	40 
    -- CP-element group 49: 	46 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (10) 
      -- CP-element group 49: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566__exit__
      -- CP-element group 49: 	 branch_block_stmt_1259/if_stmt_1567__entry__
      -- CP-element group 49: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/$exit
      -- CP-element group 49: 	 branch_block_stmt_1259/if_stmt_1567_dead_link/$entry
      -- CP-element group 49: 	 branch_block_stmt_1259/if_stmt_1567_eval_test/$entry
      -- CP-element group 49: 	 branch_block_stmt_1259/if_stmt_1567_eval_test/$exit
      -- CP-element group 49: 	 branch_block_stmt_1259/if_stmt_1567_eval_test/branch_req
      -- CP-element group 49: 	 branch_block_stmt_1259/R_cmp_1568_place
      -- CP-element group 49: 	 branch_block_stmt_1259/if_stmt_1567_if_link/$entry
      -- CP-element group 49: 	 branch_block_stmt_1259/if_stmt_1567_else_link/$entry
      -- 
    branch_req_4614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(49), ack => if_stmt_1567_branch_req_0); -- 
    convTransposeA_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(32) & convTransposeA_CP_3784_elements(40) & convTransposeA_CP_3784_elements(46) & convTransposeA_CP_3784_elements(48);
      gj_convTransposeA_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	76 
    -- CP-element group 50: 	77 
    -- CP-element group 50:  members (24) 
      -- CP-element group 50: 	 branch_block_stmt_1259/merge_stmt_1573__exit__
      -- CP-element group 50: 	 branch_block_stmt_1259/assign_stmt_1579__entry__
      -- CP-element group 50: 	 branch_block_stmt_1259/assign_stmt_1579__exit__
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody
      -- CP-element group 50: 	 branch_block_stmt_1259/if_stmt_1567_if_link/$exit
      -- CP-element group 50: 	 branch_block_stmt_1259/if_stmt_1567_if_link/if_choice_transition
      -- CP-element group 50: 	 branch_block_stmt_1259/whilex_xbody_ifx_xthen
      -- CP-element group 50: 	 branch_block_stmt_1259/assign_stmt_1579/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/assign_stmt_1579/$exit
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/Update/cr
      -- CP-element group 50: 	 branch_block_stmt_1259/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 50: 	 branch_block_stmt_1259/merge_stmt_1573_PhiReqMerge
      -- CP-element group 50: 	 branch_block_stmt_1259/merge_stmt_1573_PhiAck/$entry
      -- CP-element group 50: 	 branch_block_stmt_1259/merge_stmt_1573_PhiAck/$exit
      -- CP-element group 50: 	 branch_block_stmt_1259/merge_stmt_1573_PhiAck/dummy
      -- 
    if_choice_transition_4619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1567_branch_ack_1, ack => convTransposeA_CP_3784_elements(50)); -- 
    rr_4802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(50), ack => type_cast_1492_inst_req_0); -- 
    cr_4807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(50), ack => type_cast_1492_inst_req_1); -- 
    -- CP-element group 51:  fork  transition  place  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	53 
    -- CP-element group 51: 	55 
    -- CP-element group 51: 	57 
    -- CP-element group 51:  members (24) 
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621__entry__
      -- CP-element group 51: 	 branch_block_stmt_1259/merge_stmt_1581__exit__
      -- CP-element group 51: 	 branch_block_stmt_1259/merge_stmt_1581_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_1259/merge_stmt_1581_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_1259/merge_stmt_1581_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_1259/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_1259/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1259/merge_stmt_1581_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_1259/if_stmt_1567_else_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_1259/if_stmt_1567_else_link/else_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_1259/whilex_xbody_ifx_xelse
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/$entry
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_Update/cr
      -- 
    else_choice_transition_4623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1567_branch_ack_0, ack => convTransposeA_CP_3784_elements(51)); -- 
    rr_4639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(51), ack => type_cast_1590_inst_req_0); -- 
    cr_4644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(51), ack => type_cast_1590_inst_req_1); -- 
    cr_4658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(51), ack => type_cast_1599_inst_req_1); -- 
    cr_4672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(51), ack => type_cast_1615_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_Sample/ra
      -- 
    ra_4640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1590_inst_ack_0, ack => convTransposeA_CP_3784_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1590_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_Sample/rr
      -- 
    ca_4645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1590_inst_ack_1, ack => convTransposeA_CP_3784_elements(53)); -- 
    rr_4653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(53), ack => type_cast_1599_inst_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_Sample/ra
      -- 
    ra_4654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1599_inst_ack_0, ack => convTransposeA_CP_3784_elements(54)); -- 
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	51 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1599_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_Sample/rr
      -- 
    ca_4659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1599_inst_ack_1, ack => convTransposeA_CP_3784_elements(55)); -- 
    rr_4667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(55), ack => type_cast_1615_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_Sample/ra
      -- 
    ra_4668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1615_inst_ack_0, ack => convTransposeA_CP_3784_elements(56)); -- 
    -- CP-element group 57:  branch  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	51 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (13) 
      -- CP-element group 57: 	 branch_block_stmt_1259/if_stmt_1622__entry__
      -- CP-element group 57: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621__exit__
      -- CP-element group 57: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/$exit
      -- CP-element group 57: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1259/assign_stmt_1587_to_assign_stmt_1621/type_cast_1615_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_1259/if_stmt_1622_dead_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1259/if_stmt_1622_eval_test/$entry
      -- CP-element group 57: 	 branch_block_stmt_1259/if_stmt_1622_eval_test/$exit
      -- CP-element group 57: 	 branch_block_stmt_1259/if_stmt_1622_eval_test/branch_req
      -- CP-element group 57: 	 branch_block_stmt_1259/R_cmp86_1623_place
      -- CP-element group 57: 	 branch_block_stmt_1259/if_stmt_1622_if_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1259/if_stmt_1622_else_link/$entry
      -- 
    ca_4673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1615_inst_ack_1, ack => convTransposeA_CP_3784_elements(57)); -- 
    branch_req_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(57), ack => if_stmt_1622_branch_req_0); -- 
    -- CP-element group 58:  merge  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (15) 
      -- CP-element group 58: 	 branch_block_stmt_1259/merge_stmt_1628__exit__
      -- CP-element group 58: 	 branch_block_stmt_1259/assign_stmt_1632__entry__
      -- CP-element group 58: 	 branch_block_stmt_1259/merge_stmt_1628_PhiAck/dummy
      -- CP-element group 58: 	 branch_block_stmt_1259/merge_stmt_1628_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1259/merge_stmt_1628_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1259/merge_stmt_1628_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1259/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1259/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1259/if_stmt_1622_if_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1259/if_stmt_1622_if_link/if_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1259/ifx_xelse_whilex_xend
      -- CP-element group 58: 	 branch_block_stmt_1259/assign_stmt_1632/$entry
      -- CP-element group 58: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_Sample/req
      -- 
    if_choice_transition_4686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1622_branch_ack_1, ack => convTransposeA_CP_3784_elements(58)); -- 
    req_4703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(58), ack => WPIPE_Block0_done_1630_inst_req_0); -- 
    -- CP-element group 59:  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	65 
    -- CP-element group 59: 	66 
    -- CP-element group 59: 	68 
    -- CP-element group 59: 	69 
    -- CP-element group 59:  members (20) 
      -- CP-element group 59: 	 branch_block_stmt_1259/if_stmt_1622_else_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1259/if_stmt_1622_else_link/else_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1622_branch_ack_0, ack => convTransposeA_CP_3784_elements(59)); -- 
    rr_4747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(59), ack => type_cast_1425_inst_req_0); -- 
    cr_4752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(59), ack => type_cast_1425_inst_req_1); -- 
    rr_4770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(59), ack => type_cast_1432_inst_req_0); -- 
    cr_4775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(59), ack => type_cast_1432_inst_req_1); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_Sample/ack
      -- CP-element group 60: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_Update/req
      -- 
    ack_4704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1630_inst_ack_0, ack => convTransposeA_CP_3784_elements(60)); -- 
    req_4708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(60), ack => WPIPE_Block0_done_1630_inst_req_1); -- 
    -- CP-element group 61:  transition  place  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (16) 
      -- CP-element group 61: 	 branch_block_stmt_1259/branch_block_stmt_1259__exit__
      -- CP-element group 61: 	 branch_block_stmt_1259/assign_stmt_1632__exit__
      -- CP-element group 61: 	 branch_block_stmt_1259/return__
      -- CP-element group 61: 	 branch_block_stmt_1259/merge_stmt_1634__exit__
      -- CP-element group 61: 	 branch_block_stmt_1259/$exit
      -- CP-element group 61: 	 $exit
      -- CP-element group 61: 	 branch_block_stmt_1259/merge_stmt_1634_PhiAck/dummy
      -- CP-element group 61: 	 branch_block_stmt_1259/merge_stmt_1634_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_1259/merge_stmt_1634_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_1259/return___PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_1259/return___PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_1259/merge_stmt_1634_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_1259/assign_stmt_1632/$exit
      -- CP-element group 61: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1259/assign_stmt_1632/WPIPE_Block0_done_1630_Update/ack
      -- 
    ack_4709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1630_inst_ack_1, ack => convTransposeA_CP_3784_elements(61)); -- 
    -- CP-element group 62:  transition  output  delay-element  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	29 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/$exit
      -- CP-element group 62: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/$exit
      -- CP-element group 62: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1423_konst_delay_trans
      -- CP-element group 62: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_req
      -- 
    phi_stmt_1419_req_4720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1419_req_4720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(62), ack => phi_stmt_1419_req_0); -- 
    -- Element group convTransposeA_CP_3784_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => convTransposeA_CP_3784_elements(29), ack => convTransposeA_CP_3784_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  transition  output  delay-element  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	29 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/$exit
      -- CP-element group 63: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/$exit
      -- CP-element group 63: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1430_konst_delay_trans
      -- CP-element group 63: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_req
      -- 
    phi_stmt_1426_req_4728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1426_req_4728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(63), ack => phi_stmt_1426_req_0); -- 
    -- Element group convTransposeA_CP_3784_elements(63) is a control-delay.
    cp_element_63_delay: control_delay_element  generic map(name => " 63_delay", delay_value => 1)  port map(req => convTransposeA_CP_3784_elements(29), ack => convTransposeA_CP_3784_elements(63), clk => clk, reset =>reset);
    -- CP-element group 64:  join  transition  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	72 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1259/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(62) & convTransposeA_CP_3784_elements(63);
      gj_convTransposeA_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	59 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/Sample/ra
      -- 
    ra_4748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_0, ack => convTransposeA_CP_3784_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	59 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/Update/ca
      -- 
    ca_4753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1425_inst_ack_1, ack => convTransposeA_CP_3784_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (5) 
      -- CP-element group 67: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/$exit
      -- CP-element group 67: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/$exit
      -- CP-element group 67: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/$exit
      -- CP-element group 67: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_sources/type_cast_1425/SplitProtocol/$exit
      -- CP-element group 67: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1419/phi_stmt_1419_req
      -- 
    phi_stmt_1419_req_4754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1419_req_4754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(67), ack => phi_stmt_1419_req_1); -- 
    convTransposeA_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(65) & convTransposeA_CP_3784_elements(66);
      gj_convTransposeA_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	59 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/Sample/ra
      -- 
    ra_4771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1432_inst_ack_0, ack => convTransposeA_CP_3784_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	59 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/Update/ca
      -- 
    ca_4776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1432_inst_ack_1, ack => convTransposeA_CP_3784_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (5) 
      -- CP-element group 70: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/$exit
      -- CP-element group 70: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/$exit
      -- CP-element group 70: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_sources/type_cast_1432/SplitProtocol/$exit
      -- CP-element group 70: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1426/phi_stmt_1426_req
      -- 
    phi_stmt_1426_req_4777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1426_req_4777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(70), ack => phi_stmt_1426_req_1); -- 
    convTransposeA_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(68) & convTransposeA_CP_3784_elements(69);
      gj_convTransposeA_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1259/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(67) & convTransposeA_CP_3784_elements(70);
      gj_convTransposeA_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  merge  fork  transition  place  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	64 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1259/merge_stmt_1418_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1259/merge_stmt_1418_PhiAck/$entry
      -- 
    convTransposeA_CP_3784_elements(72) <= OrReduce(convTransposeA_CP_3784_elements(64) & convTransposeA_CP_3784_elements(71));
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1259/merge_stmt_1418_PhiAck/phi_stmt_1419_ack
      -- 
    phi_stmt_1419_ack_4782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1419_ack_0, ack => convTransposeA_CP_3784_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1259/merge_stmt_1418_PhiAck/phi_stmt_1426_ack
      -- 
    phi_stmt_1426_ack_4783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1426_ack_0, ack => convTransposeA_CP_3784_elements(74)); -- 
    -- CP-element group 75:  join  transition  place  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (10) 
      -- CP-element group 75: 	 branch_block_stmt_1259/assign_stmt_1438_to_assign_stmt_1483__exit__
      -- CP-element group 75: 	 branch_block_stmt_1259/assign_stmt_1438_to_assign_stmt_1483__entry__
      -- CP-element group 75: 	 branch_block_stmt_1259/merge_stmt_1418__exit__
      -- CP-element group 75: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 75: 	 branch_block_stmt_1259/assign_stmt_1438_to_assign_stmt_1483/$entry
      -- CP-element group 75: 	 branch_block_stmt_1259/assign_stmt_1438_to_assign_stmt_1483/$exit
      -- CP-element group 75: 	 branch_block_stmt_1259/merge_stmt_1418_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1486/$entry
      -- CP-element group 75: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/$entry
      -- 
    convTransposeA_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(73) & convTransposeA_CP_3784_elements(74);
      gj_convTransposeA_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	50 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/Sample/ra
      -- 
    ra_4803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1492_inst_ack_0, ack => convTransposeA_CP_3784_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	50 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/Update/ca
      -- 
    ca_4808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1492_inst_ack_1, ack => convTransposeA_CP_3784_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/$exit
      -- CP-element group 78: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/$exit
      -- CP-element group 78: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1492/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_1259/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_req
      -- 
    phi_stmt_1486_req_4809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1486_req_4809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(78), ack => phi_stmt_1486_req_1); -- 
    convTransposeA_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3784_elements(76) & convTransposeA_CP_3784_elements(77);
      gj_convTransposeA_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3784_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 79: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1486/$exit
      -- CP-element group 79: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_sources/type_cast_1490_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1259/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1486/phi_stmt_1486_req
      -- 
    phi_stmt_1486_req_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1486_req_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(79), ack => phi_stmt_1486_req_0); -- 
    -- Element group convTransposeA_CP_3784_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3784_elements(75), ack => convTransposeA_CP_3784_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  merge  transition  place  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1259/merge_stmt_1485_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_1259/merge_stmt_1485_PhiAck/$entry
      -- 
    convTransposeA_CP_3784_elements(80) <= OrReduce(convTransposeA_CP_3784_elements(78) & convTransposeA_CP_3784_elements(79));
    -- CP-element group 81:  fork  transition  place  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	30 
    -- CP-element group 81: 	31 
    -- CP-element group 81: 	33 
    -- CP-element group 81: 	35 
    -- CP-element group 81: 	37 
    -- CP-element group 81: 	38 
    -- CP-element group 81: 	39 
    -- CP-element group 81: 	41 
    -- CP-element group 81: 	43 
    -- CP-element group 81: 	46 
    -- CP-element group 81: 	47 
    -- CP-element group 81: 	48 
    -- CP-element group 81:  members (45) 
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566__entry__
      -- CP-element group 81: 	 branch_block_stmt_1259/merge_stmt_1485__exit__
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1512_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_update_start
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1524_final_index_sum_regn_Update/req
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1525_complete/req
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1529_Update/word_access_complete/word_0/cr
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1533_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_update_start
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/array_obj_ref_1545_final_index_sum_regn_Update/req
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/addr_of_1546_complete/req
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/ptr_deref_1549_Update/word_access_complete/word_0/cr
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1259/assign_stmt_1499_to_assign_stmt_1566/type_cast_1554_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_1259/merge_stmt_1485_PhiAck/$exit
      -- CP-element group 81: 	 branch_block_stmt_1259/merge_stmt_1485_PhiAck/phi_stmt_1486_ack
      -- 
    phi_stmt_1486_ack_4825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1486_ack_0, ack => convTransposeA_CP_3784_elements(81)); -- 
    rr_4380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => type_cast_1512_inst_req_0); -- 
    cr_4385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => type_cast_1512_inst_req_1); -- 
    req_4416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => array_obj_ref_1524_index_offset_req_1); -- 
    req_4431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => addr_of_1525_final_reg_req_1); -- 
    cr_4476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => ptr_deref_1529_load_0_req_1); -- 
    rr_4490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => type_cast_1533_inst_req_0); -- 
    cr_4495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => type_cast_1533_inst_req_1); -- 
    req_4526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => array_obj_ref_1545_index_offset_req_1); -- 
    req_4541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => addr_of_1546_final_reg_req_1); -- 
    cr_4591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => ptr_deref_1549_store_0_req_1); -- 
    rr_4600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => type_cast_1554_inst_req_0); -- 
    cr_4605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3784_elements(81), ack => type_cast_1554_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_padding_1311_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1311_word_address_0 : std_logic_vector(0 downto 0);
    signal R_shr100_1523_resized : std_logic_vector(13 downto 0);
    signal R_shr100_1523_scaled : std_logic_vector(13 downto 0);
    signal R_shr57102_1544_resized : std_logic_vector(13 downto 0);
    signal R_shr57102_1544_scaled : std_logic_vector(13 downto 0);
    signal add10_1504 : std_logic_vector(15 downto 0);
    signal add50_1509 : std_logic_vector(15 downto 0);
    signal add63_1561 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1524_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1524_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1545_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1545_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1545_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1545_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1545_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1545_root_address : std_logic_vector(13 downto 0);
    signal arrayidx59_1547 : std_logic_vector(31 downto 0);
    signal arrayidx_1526 : std_logic_vector(31 downto 0);
    signal call_1262 : std_logic_vector(15 downto 0);
    signal cmp76_1596 : std_logic_vector(0 downto 0);
    signal cmp86_1621 : std_logic_vector(0 downto 0);
    signal cmp_1566 : std_logic_vector(0 downto 0);
    signal conv53_1513 : std_logic_vector(63 downto 0);
    signal conv56_1534 : std_logic_vector(63 downto 0);
    signal conv62_1555 : std_logic_vector(31 downto 0);
    signal conv65_1362 : std_logic_vector(31 downto 0);
    signal conv73_1591 : std_logic_vector(31 downto 0);
    signal conv75_1366 : std_logic_vector(31 downto 0);
    signal conv82_1616 : std_logic_vector(31 downto 0);
    signal conv84_1388 : std_logic_vector(31 downto 0);
    signal div85_1394 : std_logic_vector(31 downto 0);
    signal div_1372 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1380 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1271 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1283 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1293 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1305 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1318 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1330 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1342 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1354 : std_logic_vector(31 downto 0);
    signal inc80_1600 : std_logic_vector(15 downto 0);
    signal inc80x_xinput_dim0x_x2_1605 : std_logic_vector(15 downto 0);
    signal inc_1587 : std_logic_vector(15 downto 0);
    signal indvar_1486 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1579 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1426 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1419 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1612 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1499 : std_logic_vector(15 downto 0);
    signal ptr_deref_1274_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1274_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1274_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1274_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1274_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1286_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1286_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1286_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1286_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1286_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1296_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1296_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1296_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1296_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1296_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1308_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1308_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1308_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1308_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1308_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1321_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1321_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1321_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1321_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1321_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1333_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1333_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1333_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1333_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1333_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1345_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1345_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1345_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1345_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1345_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1357_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1357_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1357_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1357_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1357_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1383_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1383_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1383_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1383_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1383_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1529_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1529_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1529_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1529_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1529_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1549_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1549_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1549_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1549_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1549_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1549_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr100_1519 : std_logic_vector(63 downto 0);
    signal shr57102_1540 : std_logic_vector(63 downto 0);
    signal tmp10_1473 : std_logic_vector(15 downto 0);
    signal tmp115_1438 : std_logic_vector(15 downto 0);
    signal tmp116_1443 : std_logic_vector(15 downto 0);
    signal tmp117_1448 : std_logic_vector(15 downto 0);
    signal tmp11_1478 : std_logic_vector(15 downto 0);
    signal tmp12_1483 : std_logic_vector(15 downto 0);
    signal tmp14_1297 : std_logic_vector(15 downto 0);
    signal tmp17_1309 : std_logic_vector(15 downto 0);
    signal tmp1_1275 : std_logic_vector(15 downto 0);
    signal tmp20_1312 : std_logic_vector(15 downto 0);
    signal tmp26_1322 : std_logic_vector(15 downto 0);
    signal tmp29_1334 : std_logic_vector(15 downto 0);
    signal tmp2_1405 : std_logic_vector(15 downto 0);
    signal tmp39_1346 : std_logic_vector(15 downto 0);
    signal tmp3_1453 : std_logic_vector(15 downto 0);
    signal tmp43_1358 : std_logic_vector(15 downto 0);
    signal tmp4_1458 : std_logic_vector(15 downto 0);
    signal tmp54_1530 : std_logic_vector(63 downto 0);
    signal tmp5_1287 : std_logic_vector(15 downto 0);
    signal tmp6_1411 : std_logic_vector(15 downto 0);
    signal tmp7_1416 : std_logic_vector(15 downto 0);
    signal tmp83_1384 : std_logic_vector(15 downto 0);
    signal tmp8_1463 : std_logic_vector(15 downto 0);
    signal tmp9_1468 : std_logic_vector(15 downto 0);
    signal tmp_1400 : std_logic_vector(15 downto 0);
    signal type_cast_1370_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1392_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1398_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1409_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1423_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1425_wire : std_logic_vector(15 downto 0);
    signal type_cast_1430_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1432_wire : std_logic_vector(15 downto 0);
    signal type_cast_1490_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1492_wire : std_logic_vector(15 downto 0);
    signal type_cast_1497_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1517_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1538_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1559_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1577_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1585_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1609_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_padding_1311_word_address_0 <= "0";
    array_obj_ref_1524_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1524_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1524_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1524_resized_base_address <= "00000000000000";
    array_obj_ref_1545_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1545_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1545_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1545_resized_base_address <= "00000000000000";
    iNsTr_10_1380 <= "00000000000000000000000000000011";
    iNsTr_2_1271 <= "00000000000000000000000000000101";
    iNsTr_3_1283 <= "00000000000000000000000000000100";
    iNsTr_4_1293 <= "00000000000000000000000000000000";
    iNsTr_5_1305 <= "00000000000000000000000000000100";
    iNsTr_6_1318 <= "00000000000000000000000000000001";
    iNsTr_7_1330 <= "00000000000000000000000000000101";
    iNsTr_8_1342 <= "00000000000000000000000000000101";
    iNsTr_9_1354 <= "00000000000000000000000000000100";
    ptr_deref_1274_word_offset_0 <= "0000000";
    ptr_deref_1286_word_offset_0 <= "0000000";
    ptr_deref_1296_word_offset_0 <= "0";
    ptr_deref_1308_word_offset_0 <= "0000000";
    ptr_deref_1321_word_offset_0 <= "0";
    ptr_deref_1333_word_offset_0 <= "0000000";
    ptr_deref_1345_word_offset_0 <= "0000000";
    ptr_deref_1357_word_offset_0 <= "0000000";
    ptr_deref_1383_word_offset_0 <= "0000000";
    ptr_deref_1529_word_offset_0 <= "00000000000000";
    ptr_deref_1549_word_offset_0 <= "00000000000000";
    type_cast_1370_wire_constant <= "00000000000000000000000000000001";
    type_cast_1392_wire_constant <= "00000000000000000000000000000001";
    type_cast_1398_wire_constant <= "1111111111111111";
    type_cast_1409_wire_constant <= "1111111111111111";
    type_cast_1423_wire_constant <= "0000000000000000";
    type_cast_1430_wire_constant <= "0000000000000000";
    type_cast_1490_wire_constant <= "0000000000000000";
    type_cast_1497_wire_constant <= "0000000000000100";
    type_cast_1517_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1538_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1559_wire_constant <= "00000000000000000000000000000100";
    type_cast_1577_wire_constant <= "0000000000000001";
    type_cast_1585_wire_constant <= "0000000000000001";
    type_cast_1609_wire_constant <= "0000000000000000";
    phi_stmt_1419: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1423_wire_constant & type_cast_1425_wire;
      req <= phi_stmt_1419_req_0 & phi_stmt_1419_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1419",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1419_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1419,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1419
    phi_stmt_1426: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1430_wire_constant & type_cast_1432_wire;
      req <= phi_stmt_1426_req_0 & phi_stmt_1426_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1426",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1426_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1426,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1426
    phi_stmt_1486: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1490_wire_constant & type_cast_1492_wire;
      req <= phi_stmt_1486_req_0 & phi_stmt_1486_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1486",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1486_ack_0,
          idata => idata,
          odata => indvar_1486,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1486
    -- flow-through select operator MUX_1611_inst
    input_dim1x_x2_1612 <= type_cast_1609_wire_constant when (cmp76_1596(0) /=  '0') else inc_1587;
    addr_of_1525_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1525_final_reg_req_0;
      addr_of_1525_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1525_final_reg_req_1;
      addr_of_1525_final_reg_ack_1<= rack(0);
      addr_of_1525_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1525_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1524_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1546_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1546_final_reg_req_0;
      addr_of_1546_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1546_final_reg_req_1;
      addr_of_1546_final_reg_ack_1<= rack(0);
      addr_of_1546_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1546_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1545_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx59_1547,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1361_inst_req_0;
      type_cast_1361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1361_inst_req_1;
      type_cast_1361_inst_ack_1<= rack(0);
      type_cast_1361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_1275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_1362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1365_inst_req_0;
      type_cast_1365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1365_inst_req_1;
      type_cast_1365_inst_ack_1<= rack(0);
      type_cast_1365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp5_1287,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_1366,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1387_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1387_inst_req_0;
      type_cast_1387_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1387_inst_req_1;
      type_cast_1387_inst_ack_1<= rack(0);
      type_cast_1387_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1387_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp83_1384,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_1388,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1425_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1425_inst_req_0;
      type_cast_1425_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1425_inst_req_1;
      type_cast_1425_inst_ack_1<= rack(0);
      type_cast_1425_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1425_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1425_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1432_inst_req_0;
      type_cast_1432_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1432_inst_req_1;
      type_cast_1432_inst_ack_1<= rack(0);
      type_cast_1432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc80x_xinput_dim0x_x2_1605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1432_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1492_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1492_inst_req_0;
      type_cast_1492_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1492_inst_req_1;
      type_cast_1492_inst_ack_1<= rack(0);
      type_cast_1492_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1492_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1579,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1492_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1512_inst_req_0;
      type_cast_1512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1512_inst_req_1;
      type_cast_1512_inst_ack_1<= rack(0);
      type_cast_1512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1512_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add10_1504,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1513,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1533_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1533_inst_req_0;
      type_cast_1533_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1533_inst_req_1;
      type_cast_1533_inst_ack_1<= rack(0);
      type_cast_1533_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1533_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add50_1509,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1534,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1554_inst_req_0;
      type_cast_1554_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1554_inst_req_1;
      type_cast_1554_inst_ack_1<= rack(0);
      type_cast_1554_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1499,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_1555,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1590_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1590_inst_req_0;
      type_cast_1590_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1590_inst_req_1;
      type_cast_1590_inst_ack_1<= rack(0);
      type_cast_1590_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1590_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1599_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1599_inst_req_0;
      type_cast_1599_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1599_inst_req_1;
      type_cast_1599_inst_ack_1<= rack(0);
      type_cast_1599_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1599_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp76_1596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc80_1600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1615_inst_req_0;
      type_cast_1615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1615_inst_req_1;
      type_cast_1615_inst_ack_1<= rack(0);
      type_cast_1615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc80x_xinput_dim0x_x2_1605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_1616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1311_gather_scatter
    process(LOAD_padding_1311_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1311_data_0;
      ov(15 downto 0) := iv;
      tmp20_1312 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1524_index_1_rename
    process(R_shr100_1523_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr100_1523_resized;
      ov(13 downto 0) := iv;
      R_shr100_1523_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1524_index_1_resize
    process(shr100_1519) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr100_1519;
      ov := iv(13 downto 0);
      R_shr100_1523_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1524_root_address_inst
    process(array_obj_ref_1524_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1524_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1524_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1545_index_1_rename
    process(R_shr57102_1544_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr57102_1544_resized;
      ov(13 downto 0) := iv;
      R_shr57102_1544_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1545_index_1_resize
    process(shr57102_1540) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr57102_1540;
      ov := iv(13 downto 0);
      R_shr57102_1544_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1545_root_address_inst
    process(array_obj_ref_1545_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1545_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1545_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1274_addr_0
    process(ptr_deref_1274_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1274_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1274_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1274_base_resize
    process(iNsTr_2_1271) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1271;
      ov := iv(6 downto 0);
      ptr_deref_1274_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1274_gather_scatter
    process(ptr_deref_1274_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1274_data_0;
      ov(15 downto 0) := iv;
      tmp1_1275 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1274_root_address_inst
    process(ptr_deref_1274_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1274_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1274_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1286_addr_0
    process(ptr_deref_1286_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1286_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1286_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1286_base_resize
    process(iNsTr_3_1283) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1283;
      ov := iv(6 downto 0);
      ptr_deref_1286_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1286_gather_scatter
    process(ptr_deref_1286_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1286_data_0;
      ov(15 downto 0) := iv;
      tmp5_1287 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1286_root_address_inst
    process(ptr_deref_1286_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1286_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1286_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1296_addr_0
    process(ptr_deref_1296_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1296_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1296_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1296_base_resize
    process(iNsTr_4_1293) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1293;
      ov := iv(0 downto 0);
      ptr_deref_1296_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1296_gather_scatter
    process(ptr_deref_1296_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1296_data_0;
      ov(15 downto 0) := iv;
      tmp14_1297 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1296_root_address_inst
    process(ptr_deref_1296_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1296_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1296_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1308_addr_0
    process(ptr_deref_1308_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1308_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1308_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1308_base_resize
    process(iNsTr_5_1305) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1305;
      ov := iv(6 downto 0);
      ptr_deref_1308_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1308_gather_scatter
    process(ptr_deref_1308_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1308_data_0;
      ov(15 downto 0) := iv;
      tmp17_1309 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1308_root_address_inst
    process(ptr_deref_1308_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1308_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1308_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1321_addr_0
    process(ptr_deref_1321_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1321_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1321_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1321_base_resize
    process(iNsTr_6_1318) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1318;
      ov := iv(0 downto 0);
      ptr_deref_1321_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1321_gather_scatter
    process(ptr_deref_1321_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1321_data_0;
      ov(15 downto 0) := iv;
      tmp26_1322 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1321_root_address_inst
    process(ptr_deref_1321_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1321_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1321_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1333_addr_0
    process(ptr_deref_1333_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1333_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1333_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1333_base_resize
    process(iNsTr_7_1330) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1330;
      ov := iv(6 downto 0);
      ptr_deref_1333_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1333_gather_scatter
    process(ptr_deref_1333_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1333_data_0;
      ov(15 downto 0) := iv;
      tmp29_1334 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1333_root_address_inst
    process(ptr_deref_1333_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1333_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1333_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1345_addr_0
    process(ptr_deref_1345_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1345_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1345_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1345_base_resize
    process(iNsTr_8_1342) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1342;
      ov := iv(6 downto 0);
      ptr_deref_1345_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1345_gather_scatter
    process(ptr_deref_1345_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1345_data_0;
      ov(15 downto 0) := iv;
      tmp39_1346 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1345_root_address_inst
    process(ptr_deref_1345_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1345_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1345_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1357_addr_0
    process(ptr_deref_1357_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1357_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1357_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1357_base_resize
    process(iNsTr_9_1354) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1354;
      ov := iv(6 downto 0);
      ptr_deref_1357_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1357_gather_scatter
    process(ptr_deref_1357_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1357_data_0;
      ov(15 downto 0) := iv;
      tmp43_1358 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1357_root_address_inst
    process(ptr_deref_1357_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1357_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1357_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1383_addr_0
    process(ptr_deref_1383_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1383_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1383_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1383_base_resize
    process(iNsTr_10_1380) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1380;
      ov := iv(6 downto 0);
      ptr_deref_1383_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1383_gather_scatter
    process(ptr_deref_1383_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1383_data_0;
      ov(15 downto 0) := iv;
      tmp83_1384 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1383_root_address_inst
    process(ptr_deref_1383_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1383_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1383_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1529_addr_0
    process(ptr_deref_1529_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1529_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1529_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1529_base_resize
    process(arrayidx_1526) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1526;
      ov := iv(13 downto 0);
      ptr_deref_1529_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1529_gather_scatter
    process(ptr_deref_1529_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1529_data_0;
      ov(63 downto 0) := iv;
      tmp54_1530 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1529_root_address_inst
    process(ptr_deref_1529_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1529_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1529_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1549_addr_0
    process(ptr_deref_1549_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1549_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1549_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1549_base_resize
    process(arrayidx59_1547) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx59_1547;
      ov := iv(13 downto 0);
      ptr_deref_1549_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1549_gather_scatter
    process(tmp54_1530) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp54_1530;
      ov(63 downto 0) := iv;
      ptr_deref_1549_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1549_root_address_inst
    process(ptr_deref_1549_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1549_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1549_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1567_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1566;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1567_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1567_branch_req_0,
          ack0 => if_stmt_1567_branch_ack_0,
          ack1 => if_stmt_1567_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1622_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp86_1621;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1622_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1622_branch_req_0,
          ack0 => if_stmt_1622_branch_ack_0,
          ack1 => if_stmt_1622_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1399_inst
    process(tmp29_1334) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp29_1334, type_cast_1398_wire_constant, tmp_var);
      tmp_1400 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1410_inst
    process(tmp17_1309) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp17_1309, type_cast_1409_wire_constant, tmp_var);
      tmp6_1411 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1442_inst
    process(input_dim1x_x1x_xph_1419, tmp115_1438) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1419, tmp115_1438, tmp_var);
      tmp116_1443 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1457_inst
    process(tmp2_1405, tmp3_1453) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_1405, tmp3_1453, tmp_var);
      tmp4_1458 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1467_inst
    process(tmp7_1416, tmp8_1463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp7_1416, tmp8_1463, tmp_var);
      tmp9_1468 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1477_inst
    process(tmp4_1458, tmp10_1473) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_1458, tmp10_1473, tmp_var);
      tmp11_1478 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1503_inst
    process(tmp117_1448, input_dim2x_x1_1499) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp117_1448, input_dim2x_x1_1499, tmp_var);
      add10_1504 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1508_inst
    process(tmp12_1483, input_dim2x_x1_1499) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp12_1483, input_dim2x_x1_1499, tmp_var);
      add50_1509 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1578_inst
    process(indvar_1486) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1486, type_cast_1577_wire_constant, tmp_var);
      indvarx_xnext_1579 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1586_inst
    process(input_dim1x_x1x_xph_1419) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1419, type_cast_1585_wire_constant, tmp_var);
      inc_1587 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1604_inst
    process(inc80_1600, input_dim0x_x2x_xph_1426) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc80_1600, input_dim0x_x2x_xph_1426, tmp_var);
      inc80x_xinput_dim0x_x2_1605 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1560_inst
    process(conv62_1555) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv62_1555, type_cast_1559_wire_constant, tmp_var);
      add63_1561 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1595_inst
    process(conv73_1591, div_1372) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv73_1591, div_1372, tmp_var);
      cmp76_1596 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1620_inst
    process(conv82_1616, div85_1394) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv82_1616, div85_1394, tmp_var);
      cmp86_1621 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1371_inst
    process(conv75_1366) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv75_1366, type_cast_1370_wire_constant, tmp_var);
      div_1372 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1393_inst
    process(conv84_1388) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv84_1388, type_cast_1392_wire_constant, tmp_var);
      div85_1394 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1518_inst
    process(conv53_1513) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv53_1513, type_cast_1517_wire_constant, tmp_var);
      shr100_1519 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1539_inst
    process(conv56_1534) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv56_1534, type_cast_1538_wire_constant, tmp_var);
      shr57102_1540 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1437_inst
    process(tmp5_1287, input_dim0x_x2x_xph_1426) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp5_1287, input_dim0x_x2x_xph_1426, tmp_var);
      tmp115_1438 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1447_inst
    process(tmp1_1275, tmp116_1443) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1275, tmp116_1443, tmp_var);
      tmp117_1448 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1452_inst
    process(tmp26_1322, input_dim1x_x1x_xph_1419) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp26_1322, input_dim1x_x1x_xph_1419, tmp_var);
      tmp3_1453 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1462_inst
    process(tmp14_1297, input_dim0x_x2x_xph_1426) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_1297, input_dim0x_x2x_xph_1426, tmp_var);
      tmp8_1463 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1472_inst
    process(tmp43_1358, tmp9_1468) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp43_1358, tmp9_1468, tmp_var);
      tmp10_1473 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1482_inst
    process(tmp39_1346, tmp11_1478) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp39_1346, tmp11_1478, tmp_var);
      tmp12_1483 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1498_inst
    process(indvar_1486) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1486, type_cast_1497_wire_constant, tmp_var);
      input_dim2x_x1_1499 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1404_inst
    process(tmp_1400, tmp20_1312) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp_1400, tmp20_1312, tmp_var);
      tmp2_1405 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1415_inst
    process(tmp6_1411, tmp20_1312) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp6_1411, tmp20_1312, tmp_var);
      tmp7_1416 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1565_inst
    process(add63_1561, conv65_1362) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add63_1561, conv65_1362, tmp_var);
      cmp_1566 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1524_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr100_1523_scaled;
      array_obj_ref_1524_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1524_index_offset_req_0;
      array_obj_ref_1524_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1524_index_offset_req_1;
      array_obj_ref_1524_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1545_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr57102_1544_scaled;
      array_obj_ref_1545_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1545_index_offset_req_0;
      array_obj_ref_1545_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1545_index_offset_req_1;
      array_obj_ref_1545_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : LOAD_padding_1311_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1311_load_0_req_0;
      LOAD_padding_1311_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1311_load_0_req_1;
      LOAD_padding_1311_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1311_word_address_0;
      LOAD_padding_1311_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1286_load_0 ptr_deref_1383_load_0 ptr_deref_1274_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1286_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1383_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1274_load_0_req_0;
      ptr_deref_1286_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1383_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1274_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1286_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1383_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1274_load_0_req_1;
      ptr_deref_1286_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1383_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1274_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1286_word_address_0 & ptr_deref_1383_word_address_0 & ptr_deref_1274_word_address_0;
      ptr_deref_1286_data_0 <= data_out(47 downto 32);
      ptr_deref_1383_data_0 <= data_out(31 downto 16);
      ptr_deref_1274_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1296_load_0 ptr_deref_1321_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1296_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1321_load_0_req_0;
      ptr_deref_1296_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1321_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1296_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1321_load_0_req_1;
      ptr_deref_1296_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1321_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1296_word_address_0 & ptr_deref_1321_word_address_0;
      ptr_deref_1296_data_0 <= data_out(31 downto 16);
      ptr_deref_1321_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1308_load_0 ptr_deref_1333_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1308_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1333_load_0_req_0;
      ptr_deref_1308_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1333_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1308_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1333_load_0_req_1;
      ptr_deref_1308_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1333_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1308_word_address_0 & ptr_deref_1333_word_address_0;
      ptr_deref_1308_data_0 <= data_out(31 downto 16);
      ptr_deref_1333_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1345_load_0 ptr_deref_1357_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1345_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1357_load_0_req_0;
      ptr_deref_1345_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1357_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1345_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1357_load_0_req_1;
      ptr_deref_1345_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1357_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1345_word_address_0 & ptr_deref_1357_word_address_0;
      ptr_deref_1345_data_0 <= data_out(31 downto 16);
      ptr_deref_1357_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1529_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1529_load_0_req_0;
      ptr_deref_1529_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1529_load_0_req_1;
      ptr_deref_1529_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1529_word_address_0;
      ptr_deref_1529_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1549_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1549_store_0_req_0;
      ptr_deref_1549_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1549_store_0_req_1;
      ptr_deref_1549_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1549_word_address_0;
      data_in <= ptr_deref_1549_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1261_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_start_1261_inst_req_0;
      RPIPE_Block0_start_1261_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_start_1261_inst_req_1;
      RPIPE_Block0_start_1261_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1262 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1630_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1630_inst_req_0;
      WPIPE_Block0_done_1630_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1630_inst_req_1;
      WPIPE_Block0_done_1630_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1262;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4866_start: Boolean;
  signal convTransposeB_CP_4866_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1653_load_0_req_0 : boolean;
  signal ptr_deref_1681_load_0_ack_0 : boolean;
  signal type_cast_1799_inst_req_1 : boolean;
  signal ptr_deref_1653_load_0_ack_0 : boolean;
  signal ptr_deref_1671_load_0_req_1 : boolean;
  signal type_cast_1806_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1640_inst_ack_1 : boolean;
  signal ptr_deref_1681_load_0_req_1 : boolean;
  signal RPIPE_Block1_start_1640_inst_req_1 : boolean;
  signal ptr_deref_1671_load_0_ack_1 : boolean;
  signal ptr_deref_1653_load_0_ack_1 : boolean;
  signal RPIPE_Block1_start_1640_inst_req_0 : boolean;
  signal ptr_deref_1681_load_0_ack_1 : boolean;
  signal ptr_deref_1681_load_0_req_0 : boolean;
  signal RPIPE_Block1_start_1640_inst_ack_0 : boolean;
  signal ptr_deref_1671_load_0_req_0 : boolean;
  signal ptr_deref_1671_load_0_ack_0 : boolean;
  signal ptr_deref_1653_load_0_req_1 : boolean;
  signal type_cast_1799_inst_ack_1 : boolean;
  signal phi_stmt_1860_ack_0 : boolean;
  signal type_cast_1797_inst_req_0 : boolean;
  signal type_cast_1797_inst_ack_0 : boolean;
  signal type_cast_1806_inst_ack_0 : boolean;
  signal phi_stmt_1794_req_1 : boolean;
  signal ptr_deref_1693_load_0_req_0 : boolean;
  signal ptr_deref_1693_load_0_ack_0 : boolean;
  signal ptr_deref_1693_load_0_req_1 : boolean;
  signal ptr_deref_1693_load_0_ack_1 : boolean;
  signal LOAD_padding_1696_load_0_req_0 : boolean;
  signal LOAD_padding_1696_load_0_ack_0 : boolean;
  signal LOAD_padding_1696_load_0_req_1 : boolean;
  signal LOAD_padding_1696_load_0_ack_1 : boolean;
  signal ptr_deref_1706_load_0_req_0 : boolean;
  signal ptr_deref_1706_load_0_ack_0 : boolean;
  signal ptr_deref_1706_load_0_req_1 : boolean;
  signal ptr_deref_1706_load_0_ack_1 : boolean;
  signal ptr_deref_1718_load_0_req_0 : boolean;
  signal ptr_deref_1718_load_0_ack_0 : boolean;
  signal ptr_deref_1718_load_0_req_1 : boolean;
  signal ptr_deref_1718_load_0_ack_1 : boolean;
  signal ptr_deref_1730_load_0_req_0 : boolean;
  signal ptr_deref_1730_load_0_ack_0 : boolean;
  signal ptr_deref_1730_load_0_req_1 : boolean;
  signal ptr_deref_1730_load_0_ack_1 : boolean;
  signal ptr_deref_1742_load_0_req_0 : boolean;
  signal ptr_deref_1742_load_0_ack_0 : boolean;
  signal ptr_deref_1742_load_0_req_1 : boolean;
  signal ptr_deref_1742_load_0_ack_1 : boolean;
  signal type_cast_1746_inst_req_0 : boolean;
  signal type_cast_1746_inst_ack_0 : boolean;
  signal type_cast_1746_inst_req_1 : boolean;
  signal type_cast_1746_inst_ack_1 : boolean;
  signal ptr_deref_1758_load_0_req_0 : boolean;
  signal ptr_deref_1758_load_0_ack_0 : boolean;
  signal ptr_deref_1758_load_0_req_1 : boolean;
  signal ptr_deref_1758_load_0_ack_1 : boolean;
  signal type_cast_1762_inst_req_0 : boolean;
  signal type_cast_1762_inst_ack_0 : boolean;
  signal type_cast_1762_inst_req_1 : boolean;
  signal type_cast_1762_inst_ack_1 : boolean;
  signal phi_stmt_1860_req_1 : boolean;
  signal type_cast_1886_inst_req_0 : boolean;
  signal type_cast_1886_inst_ack_0 : boolean;
  signal type_cast_1886_inst_req_1 : boolean;
  signal type_cast_1886_inst_ack_1 : boolean;
  signal array_obj_ref_1898_index_offset_req_0 : boolean;
  signal array_obj_ref_1898_index_offset_ack_0 : boolean;
  signal array_obj_ref_1898_index_offset_req_1 : boolean;
  signal array_obj_ref_1898_index_offset_ack_1 : boolean;
  signal phi_stmt_1860_req_0 : boolean;
  signal addr_of_1899_final_reg_req_0 : boolean;
  signal addr_of_1899_final_reg_ack_0 : boolean;
  signal addr_of_1899_final_reg_req_1 : boolean;
  signal addr_of_1899_final_reg_ack_1 : boolean;
  signal type_cast_1863_inst_ack_1 : boolean;
  signal ptr_deref_1903_load_0_req_0 : boolean;
  signal type_cast_1863_inst_req_1 : boolean;
  signal ptr_deref_1903_load_0_ack_0 : boolean;
  signal type_cast_1799_inst_ack_0 : boolean;
  signal ptr_deref_1903_load_0_req_1 : boolean;
  signal ptr_deref_1903_load_0_ack_1 : boolean;
  signal type_cast_1863_inst_ack_0 : boolean;
  signal type_cast_1907_inst_req_0 : boolean;
  signal type_cast_1907_inst_ack_0 : boolean;
  signal type_cast_1907_inst_req_1 : boolean;
  signal type_cast_1907_inst_ack_1 : boolean;
  signal type_cast_1863_inst_req_0 : boolean;
  signal array_obj_ref_1919_index_offset_req_0 : boolean;
  signal array_obj_ref_1919_index_offset_ack_0 : boolean;
  signal array_obj_ref_1919_index_offset_req_1 : boolean;
  signal array_obj_ref_1919_index_offset_ack_1 : boolean;
  signal phi_stmt_1800_req_1 : boolean;
  signal addr_of_1920_final_reg_req_0 : boolean;
  signal addr_of_1920_final_reg_ack_0 : boolean;
  signal addr_of_1920_final_reg_req_1 : boolean;
  signal addr_of_1920_final_reg_ack_1 : boolean;
  signal type_cast_1799_inst_req_0 : boolean;
  signal ptr_deref_1923_store_0_req_0 : boolean;
  signal ptr_deref_1923_store_0_ack_0 : boolean;
  signal ptr_deref_1923_store_0_req_1 : boolean;
  signal ptr_deref_1923_store_0_ack_1 : boolean;
  signal phi_stmt_1800_ack_0 : boolean;
  signal type_cast_1928_inst_req_0 : boolean;
  signal type_cast_1928_inst_ack_0 : boolean;
  signal type_cast_1928_inst_req_1 : boolean;
  signal type_cast_1928_inst_ack_1 : boolean;
  signal phi_stmt_1794_ack_0 : boolean;
  signal if_stmt_1941_branch_req_0 : boolean;
  signal phi_stmt_1794_req_0 : boolean;
  signal if_stmt_1941_branch_ack_1 : boolean;
  signal type_cast_1797_inst_ack_1 : boolean;
  signal if_stmt_1941_branch_ack_0 : boolean;
  signal type_cast_1797_inst_req_1 : boolean;
  signal type_cast_1993_inst_req_0 : boolean;
  signal type_cast_1993_inst_ack_0 : boolean;
  signal type_cast_1993_inst_req_1 : boolean;
  signal type_cast_1993_inst_ack_1 : boolean;
  signal type_cast_1806_inst_ack_1 : boolean;
  signal type_cast_1806_inst_req_1 : boolean;
  signal if_stmt_2000_branch_req_0 : boolean;
  signal if_stmt_2000_branch_ack_1 : boolean;
  signal if_stmt_2000_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2008_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2008_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2008_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2008_inst_ack_1 : boolean;
  signal phi_stmt_1800_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4866_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4866_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4866_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4866_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4866: Block -- control-path 
    signal convTransposeB_CP_4866_elements: BooleanArray(77 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4866_elements(0) <= convTransposeB_CP_4866_start;
    convTransposeB_CP_4866_symbol <= convTransposeB_CP_4866_elements(55);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1638/assign_stmt_1641/$entry
      -- CP-element group 0: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1638/$entry
      -- CP-element group 0: 	 branch_block_stmt_1638/branch_block_stmt_1638__entry__
      -- CP-element group 0: 	 branch_block_stmt_1638/assign_stmt_1641__entry__
      -- 
    rr_4914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(0), ack => RPIPE_Block1_start_1640_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_Update/$entry
      -- 
    ra_4915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1640_inst_ack_0, ack => convTransposeB_CP_4866_elements(1)); -- 
    cr_4919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(1), ack => RPIPE_Block1_start_1640_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2:  members (259) 
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1641/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1641/RPIPE_Block1_start_1640_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1641__exit__
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791__entry__
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_Update/cr
      -- 
    ca_4920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1640_inst_ack_1, ack => convTransposeB_CP_4866_elements(2)); -- 
    rr_4956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1653_load_0_req_0); -- 
    cr_5017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1671_load_0_req_1); -- 
    cr_5067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1681_load_0_req_1); -- 
    rr_5056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1681_load_0_req_0); -- 
    rr_5006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1671_load_0_req_0); -- 
    cr_4967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1653_load_0_req_1); -- 
    rr_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1693_load_0_req_0); -- 
    cr_5117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1693_load_0_req_1); -- 
    rr_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => LOAD_padding_1696_load_0_req_0); -- 
    cr_5150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => LOAD_padding_1696_load_0_req_1); -- 
    rr_5189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1706_load_0_req_0); -- 
    cr_5200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1706_load_0_req_1); -- 
    rr_5239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1718_load_0_req_0); -- 
    cr_5250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1718_load_0_req_1); -- 
    rr_5289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1730_load_0_req_0); -- 
    cr_5300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1730_load_0_req_1); -- 
    rr_5339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1742_load_0_req_0); -- 
    cr_5350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1742_load_0_req_1); -- 
    cr_5369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => type_cast_1746_inst_req_1); -- 
    rr_5403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1758_load_0_req_0); -- 
    cr_5414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => ptr_deref_1758_load_0_req_1); -- 
    cr_5433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(2), ack => type_cast_1762_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Sample/word_access_start/$exit
      -- 
    ra_4957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1653_load_0_ack_0, ack => convTransposeB_CP_4866_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	27 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/ptr_deref_1653_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/ptr_deref_1653_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/ptr_deref_1653_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/ptr_deref_1653_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1653_update_completed_
      -- 
    ca_4968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1653_load_0_ack_1, ack => convTransposeB_CP_4866_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Sample/word_access_start/word_0/ra
      -- 
    ra_5007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1671_load_0_ack_0, ack => convTransposeB_CP_4866_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/ptr_deref_1671_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/ptr_deref_1671_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/ptr_deref_1671_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1671_Update/ptr_deref_1671_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_Sample/rr
      -- 
    ca_5018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1671_load_0_ack_1, ack => convTransposeB_CP_4866_elements(6)); -- 
    rr_5364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(6), ack => type_cast_1746_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Sample/word_access_start/$exit
      -- 
    ra_5057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1681_load_0_ack_0, ack => convTransposeB_CP_4866_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	27 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/ptr_deref_1681_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/ptr_deref_1681_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/ptr_deref_1681_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1681_Update/ptr_deref_1681_Merge/merge_ack
      -- 
    ca_5068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1681_load_0_ack_1, ack => convTransposeB_CP_4866_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Sample/word_access_start/word_0/ra
      -- 
    ra_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1693_load_0_ack_0, ack => convTransposeB_CP_4866_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	27 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/ptr_deref_1693_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/ptr_deref_1693_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/ptr_deref_1693_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1693_Update/ptr_deref_1693_Merge/merge_ack
      -- 
    ca_5118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1693_load_0_ack_1, ack => convTransposeB_CP_4866_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Sample/word_access_start/word_0/ra
      -- 
    ra_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1696_load_0_ack_0, ack => convTransposeB_CP_4866_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	27 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/LOAD_padding_1696_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/LOAD_padding_1696_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/LOAD_padding_1696_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/LOAD_padding_1696_Update/LOAD_padding_1696_Merge/merge_ack
      -- 
    ca_5151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1696_load_0_ack_1, ack => convTransposeB_CP_4866_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Sample/word_access_start/word_0/ra
      -- 
    ra_5190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1706_load_0_ack_0, ack => convTransposeB_CP_4866_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	27 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/ptr_deref_1706_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/ptr_deref_1706_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/ptr_deref_1706_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1706_Update/ptr_deref_1706_Merge/merge_ack
      -- 
    ca_5201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1706_load_0_ack_1, ack => convTransposeB_CP_4866_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Sample/word_access_start/word_0/ra
      -- 
    ra_5240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1718_load_0_ack_0, ack => convTransposeB_CP_4866_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	27 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/ptr_deref_1718_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/ptr_deref_1718_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/ptr_deref_1718_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1718_Update/ptr_deref_1718_Merge/merge_ack
      -- 
    ca_5251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1718_load_0_ack_1, ack => convTransposeB_CP_4866_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Sample/word_access_start/word_0/ra
      -- 
    ra_5290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1730_load_0_ack_0, ack => convTransposeB_CP_4866_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	27 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/ptr_deref_1730_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/ptr_deref_1730_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/ptr_deref_1730_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1730_Update/ptr_deref_1730_Merge/merge_ack
      -- 
    ca_5301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1730_load_0_ack_1, ack => convTransposeB_CP_4866_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Sample/word_access_start/word_0/ra
      -- 
    ra_5340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1742_load_0_ack_0, ack => convTransposeB_CP_4866_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	27 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/ptr_deref_1742_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/ptr_deref_1742_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/ptr_deref_1742_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1742_Update/ptr_deref_1742_Merge/merge_ack
      -- 
    ca_5351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1742_load_0_ack_1, ack => convTransposeB_CP_4866_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_Sample/ra
      -- 
    ra_5365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1746_inst_ack_0, ack => convTransposeB_CP_4866_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1746_Update/ca
      -- 
    ca_5370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1746_inst_ack_1, ack => convTransposeB_CP_4866_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Sample/word_access_start/word_0/ra
      -- 
    ra_5404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1758_load_0_ack_0, ack => convTransposeB_CP_4866_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (12) 
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/ptr_deref_1758_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/ptr_deref_1758_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/ptr_deref_1758_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/ptr_deref_1758_Update/ptr_deref_1758_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_Sample/rr
      -- 
    ca_5415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1758_load_0_ack_1, ack => convTransposeB_CP_4866_elements(24)); -- 
    rr_5428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(24), ack => type_cast_1762_inst_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_Sample/ra
      -- 
    ra_5429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1762_inst_ack_0, ack => convTransposeB_CP_4866_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/type_cast_1762_Update/ca
      -- 
    ca_5434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1762_inst_ack_1, ack => convTransposeB_CP_4866_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  place  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	18 
    -- CP-element group 27: 	20 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	26 
    -- CP-element group 27: 	10 
    -- CP-element group 27: 	12 
    -- CP-element group 27: 	14 
    -- CP-element group 27: 	16 
    -- CP-element group 27: 	8 
    -- CP-element group 27: 	4 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	56 
    -- CP-element group 27: 	57 
    -- CP-element group 27: 	58 
    -- CP-element group 27:  members (14) 
      -- CP-element group 27: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791/$exit
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1638/assign_stmt_1650_to_assign_stmt_1791__exit__
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Update/cr
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/$entry
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/$entry
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/$entry
      -- CP-element group 27: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/$entry
      -- 
    rr_5776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(27), ack => type_cast_1797_inst_req_0); -- 
    cr_5781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(27), ack => type_cast_1797_inst_req_1); -- 
    convTransposeB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(18) & convTransposeB_CP_4866_elements(20) & convTransposeB_CP_4866_elements(22) & convTransposeB_CP_4866_elements(26) & convTransposeB_CP_4866_elements(10) & convTransposeB_CP_4866_elements(12) & convTransposeB_CP_4866_elements(14) & convTransposeB_CP_4866_elements(16) & convTransposeB_CP_4866_elements(8) & convTransposeB_CP_4866_elements(4);
      gj_convTransposeB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	77 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_Sample/ra
      -- 
    ra_5449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1886_inst_ack_0, ack => convTransposeB_CP_4866_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	77 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (16) 
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_resized_1
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_scaled_1
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_computed_1
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_resize_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_resize_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_resize_1/index_resize_req
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_resize_1/index_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_scale_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_scale_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_scale_1/scale_rename_req
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_index_scale_1/scale_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_Sample/req
      -- 
    ca_5454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1886_inst_ack_1, ack => convTransposeB_CP_4866_elements(29)); -- 
    req_5479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(29), ack => array_obj_ref_1898_index_offset_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	47 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_sample_complete
      -- CP-element group 30: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_Sample/ack
      -- 
    ack_5480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1898_index_offset_ack_0, ack => convTransposeB_CP_4866_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	77 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (11) 
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_offset_calculated
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_request/$entry
      -- CP-element group 31: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_request/req
      -- 
    ack_5485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1898_index_offset_ack_1, ack => convTransposeB_CP_4866_elements(31)); -- 
    req_5494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(31), ack => addr_of_1899_final_reg_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_request/$exit
      -- CP-element group 32: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_request/ack
      -- 
    ack_5495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1899_final_reg_ack_0, ack => convTransposeB_CP_4866_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	77 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (24) 
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_complete/ack
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_word_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_root_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_address_resized
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_addr_resize/$entry
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_addr_resize/$exit
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_addr_resize/base_resize_req
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_addr_resize/base_resize_ack
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_plus_offset/$entry
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_plus_offset/$exit
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_base_plus_offset/sum_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_word_addrgen/$entry
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_word_addrgen/$exit
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_word_addrgen/root_register_req
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_word_addrgen/root_register_ack
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Sample/word_access_start/$entry
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Sample/word_access_start/word_0/$entry
      -- CP-element group 33: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Sample/word_access_start/word_0/rr
      -- 
    ack_5500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1899_final_reg_ack_1, ack => convTransposeB_CP_4866_elements(33)); -- 
    rr_5533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(33), ack => ptr_deref_1903_load_0_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Sample/word_access_start/$exit
      -- CP-element group 34: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Sample/word_access_start/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Sample/word_access_start/word_0/ra
      -- 
    ra_5534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1903_load_0_ack_0, ack => convTransposeB_CP_4866_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	77 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	42 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/word_access_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/word_access_complete/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/word_access_complete/word_0/ca
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/ptr_deref_1903_Merge/$entry
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/ptr_deref_1903_Merge/$exit
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/ptr_deref_1903_Merge/merge_req
      -- CP-element group 35: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/ptr_deref_1903_Merge/merge_ack
      -- 
    ca_5545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1903_load_0_ack_1, ack => convTransposeB_CP_4866_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	77 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_Sample/ra
      -- 
    ra_5559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_0, ack => convTransposeB_CP_4866_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	77 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_resized_1
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_scaled_1
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_computed_1
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_resize_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_resize_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_resize_1/index_resize_req
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_resize_1/index_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_scale_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_scale_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_scale_1/scale_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_index_scale_1/scale_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_Sample/req
      -- 
    ca_5564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_1, ack => convTransposeB_CP_4866_elements(37)); -- 
    req_5589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(37), ack => array_obj_ref_1919_index_offset_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_sample_complete
      -- CP-element group 38: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_Sample/ack
      -- 
    ack_5590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1919_index_offset_ack_0, ack => convTransposeB_CP_4866_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	77 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (11) 
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_offset_calculated
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_request/$entry
      -- CP-element group 39: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_request/req
      -- 
    ack_5595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1919_index_offset_ack_1, ack => convTransposeB_CP_4866_elements(39)); -- 
    req_5604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(39), ack => addr_of_1920_final_reg_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_request/$exit
      -- CP-element group 40: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_request/ack
      -- 
    ack_5605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1920_final_reg_ack_0, ack => convTransposeB_CP_4866_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	77 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (19) 
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_complete/ack
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_word_addrgen/root_register_ack
      -- 
    ack_5610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1920_final_reg_ack_1, ack => convTransposeB_CP_4866_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	35 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/ptr_deref_1923_Split/$entry
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/ptr_deref_1923_Split/$exit
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/ptr_deref_1923_Split/split_req
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/ptr_deref_1923_Split/split_ack
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/word_access_start/word_0/rr
      -- 
    rr_5648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(42), ack => ptr_deref_1923_store_0_req_0); -- 
    convTransposeB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(41) & convTransposeB_CP_4866_elements(35);
      gj_convTransposeB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Sample/word_access_start/word_0/ra
      -- 
    ra_5649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1923_store_0_ack_0, ack => convTransposeB_CP_4866_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	77 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Update/word_access_complete/word_0/ca
      -- 
    ca_5660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1923_store_0_ack_1, ack => convTransposeB_CP_4866_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	77 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_Sample/ra
      -- 
    ra_5669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1928_inst_ack_0, ack => convTransposeB_CP_4866_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	77 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_Update/ca
      -- 
    ca_5674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1928_inst_ack_1, ack => convTransposeB_CP_4866_elements(46)); -- 
    -- CP-element group 47:  branch  join  transition  place  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	30 
    -- CP-element group 47: 	38 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (10) 
      -- CP-element group 47: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940__exit__
      -- CP-element group 47: 	 branch_block_stmt_1638/if_stmt_1941__entry__
      -- CP-element group 47: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/$exit
      -- CP-element group 47: 	 branch_block_stmt_1638/if_stmt_1941_dead_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_1638/if_stmt_1941_eval_test/$entry
      -- CP-element group 47: 	 branch_block_stmt_1638/if_stmt_1941_eval_test/$exit
      -- CP-element group 47: 	 branch_block_stmt_1638/if_stmt_1941_eval_test/branch_req
      -- CP-element group 47: 	 branch_block_stmt_1638/R_cmp_1942_place
      -- CP-element group 47: 	 branch_block_stmt_1638/if_stmt_1941_if_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_1638/if_stmt_1941_else_link/$entry
      -- 
    branch_req_5682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(47), ack => if_stmt_1941_branch_req_0); -- 
    convTransposeB_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(30) & convTransposeB_CP_4866_elements(38) & convTransposeB_CP_4866_elements(44) & convTransposeB_CP_4866_elements(46);
      gj_convTransposeB_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48: 	73 
    -- CP-element group 48:  members (24) 
      -- CP-element group 48: 	 branch_block_stmt_1638/assign_stmt_1953__entry__
      -- CP-element group 48: 	 branch_block_stmt_1638/assign_stmt_1953__exit__
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody
      -- CP-element group 48: 	 branch_block_stmt_1638/merge_stmt_1947__exit__
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Update/cr
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/merge_stmt_1947_PhiReqMerge
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/merge_stmt_1947_PhiAck/dummy
      -- CP-element group 48: 	 branch_block_stmt_1638/merge_stmt_1947_PhiAck/$exit
      -- CP-element group 48: 	 branch_block_stmt_1638/if_stmt_1941_if_link/$exit
      -- CP-element group 48: 	 branch_block_stmt_1638/if_stmt_1941_if_link/if_choice_transition
      -- CP-element group 48: 	 branch_block_stmt_1638/merge_stmt_1947_PhiAck/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/whilex_xbody_ifx_xthen
      -- CP-element group 48: 	 branch_block_stmt_1638/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 48: 	 branch_block_stmt_1638/assign_stmt_1953/$entry
      -- CP-element group 48: 	 branch_block_stmt_1638/assign_stmt_1953/$exit
      -- CP-element group 48: 	 branch_block_stmt_1638/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- 
    if_choice_transition_5687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1941_branch_ack_1, ack => convTransposeB_CP_4866_elements(48)); -- 
    cr_5862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(48), ack => type_cast_1863_inst_req_1); -- 
    rr_5857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(48), ack => type_cast_1863_inst_req_0); -- 
    -- CP-element group 49:  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (18) 
      -- CP-element group 49: 	 branch_block_stmt_1638/merge_stmt_1955__exit__
      -- CP-element group 49: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999__entry__
      -- CP-element group 49: 	 branch_block_stmt_1638/merge_stmt_1955_PhiReqMerge
      -- CP-element group 49: 	 branch_block_stmt_1638/merge_stmt_1955_PhiAck/dummy
      -- CP-element group 49: 	 branch_block_stmt_1638/merge_stmt_1955_PhiAck/$exit
      -- CP-element group 49: 	 branch_block_stmt_1638/merge_stmt_1955_PhiAck/$entry
      -- CP-element group 49: 	 branch_block_stmt_1638/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 49: 	 branch_block_stmt_1638/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_1638/if_stmt_1941_else_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_1638/if_stmt_1941_else_link/else_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_1638/whilex_xbody_ifx_xelse
      -- CP-element group 49: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/$entry
      -- CP-element group 49: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_Update/cr
      -- 
    else_choice_transition_5691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1941_branch_ack_0, ack => convTransposeB_CP_4866_elements(49)); -- 
    rr_5707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(49), ack => type_cast_1993_inst_req_0); -- 
    cr_5712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(49), ack => type_cast_1993_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_Sample/ra
      -- 
    ra_5708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_0, ack => convTransposeB_CP_4866_elements(50)); -- 
    -- CP-element group 51:  branch  transition  place  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_1638/if_stmt_2000__entry__
      -- CP-element group 51: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999__exit__
      -- CP-element group 51: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/$exit
      -- CP-element group 51: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1638/assign_stmt_1961_to_assign_stmt_1999/type_cast_1993_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1638/if_stmt_2000_dead_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_1638/if_stmt_2000_eval_test/$entry
      -- CP-element group 51: 	 branch_block_stmt_1638/if_stmt_2000_eval_test/$exit
      -- CP-element group 51: 	 branch_block_stmt_1638/if_stmt_2000_eval_test/branch_req
      -- CP-element group 51: 	 branch_block_stmt_1638/R_cmp100_2001_place
      -- CP-element group 51: 	 branch_block_stmt_1638/if_stmt_2000_if_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_1638/if_stmt_2000_else_link/$entry
      -- 
    ca_5713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_1, ack => convTransposeB_CP_4866_elements(51)); -- 
    branch_req_5721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(51), ack => if_stmt_2000_branch_req_0); -- 
    -- CP-element group 52:  merge  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (15) 
      -- CP-element group 52: 	 branch_block_stmt_1638/assign_stmt_2010__entry__
      -- CP-element group 52: 	 branch_block_stmt_1638/merge_stmt_2006_PhiReqMerge
      -- CP-element group 52: 	 branch_block_stmt_1638/merge_stmt_2006__exit__
      -- CP-element group 52: 	 branch_block_stmt_1638/merge_stmt_2006_PhiAck/$entry
      -- CP-element group 52: 	 branch_block_stmt_1638/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 52: 	 branch_block_stmt_1638/merge_stmt_2006_PhiAck/$exit
      -- CP-element group 52: 	 branch_block_stmt_1638/merge_stmt_2006_PhiAck/dummy
      -- CP-element group 52: 	 branch_block_stmt_1638/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_1638/if_stmt_2000_if_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_1638/if_stmt_2000_if_link/if_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_1638/ifx_xelse_whilex_xend
      -- CP-element group 52: 	 branch_block_stmt_1638/assign_stmt_2010/$entry
      -- CP-element group 52: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_Sample/req
      -- 
    if_choice_transition_5726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2000_branch_ack_1, ack => convTransposeB_CP_4866_elements(52)); -- 
    req_5743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(52), ack => WPIPE_Block1_done_2008_inst_req_0); -- 
    -- CP-element group 53:  fork  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	61 
    -- CP-element group 53: 	62 
    -- CP-element group 53: 	64 
    -- CP-element group 53: 	65 
    -- CP-element group 53:  members (20) 
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1638/if_stmt_2000_else_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_1638/if_stmt_2000_else_link/else_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter
      -- 
    else_choice_transition_5730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2000_branch_ack_0, ack => convTransposeB_CP_4866_elements(53)); -- 
    cr_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(53), ack => type_cast_1799_inst_req_1); -- 
    rr_5802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(53), ack => type_cast_1806_inst_req_0); -- 
    rr_5825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(53), ack => type_cast_1799_inst_req_0); -- 
    cr_5807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(53), ack => type_cast_1806_inst_req_1); -- 
    -- CP-element group 54:  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_Update/req
      -- 
    ack_5744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2008_inst_ack_0, ack => convTransposeB_CP_4866_elements(54)); -- 
    req_5748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(54), ack => WPIPE_Block1_done_2008_inst_req_1); -- 
    -- CP-element group 55:  transition  place  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (16) 
      -- CP-element group 55: 	 branch_block_stmt_1638/assign_stmt_2010__exit__
      -- CP-element group 55: 	 branch_block_stmt_1638/return__
      -- CP-element group 55: 	 branch_block_stmt_1638/merge_stmt_2012__exit__
      -- CP-element group 55: 	 branch_block_stmt_1638/merge_stmt_2012_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_1638/return___PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_1638/return___PhiReq/$exit
      -- CP-element group 55: 	 $exit
      -- CP-element group 55: 	 branch_block_stmt_1638/$exit
      -- CP-element group 55: 	 branch_block_stmt_1638/branch_block_stmt_1638__exit__
      -- CP-element group 55: 	 branch_block_stmt_1638/merge_stmt_2012_PhiAck/dummy
      -- CP-element group 55: 	 branch_block_stmt_1638/merge_stmt_2012_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_1638/merge_stmt_2012_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_1638/assign_stmt_2010/$exit
      -- CP-element group 55: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1638/assign_stmt_2010/WPIPE_Block1_done_2008_Update/ack
      -- 
    ack_5749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2008_inst_ack_1, ack => convTransposeB_CP_4866_elements(55)); -- 
    -- CP-element group 56:  transition  output  delay-element  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	27 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	60 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/$exit
      -- CP-element group 56: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1804_konst_delay_trans
      -- CP-element group 56: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_req
      -- 
    phi_stmt_1800_req_5760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1800_req_5760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(56), ack => phi_stmt_1800_req_0); -- 
    -- Element group convTransposeB_CP_4866_elements(56) is a control-delay.
    cp_element_56_delay: control_delay_element  generic map(name => " 56_delay", delay_value => 1)  port map(req => convTransposeB_CP_4866_elements(27), ack => convTransposeB_CP_4866_elements(56), clk => clk, reset =>reset);
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	27 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Sample/$exit
      -- 
    ra_5777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1797_inst_ack_0, ack => convTransposeB_CP_4866_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	27 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/Update/$exit
      -- 
    ca_5782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1797_inst_ack_1, ack => convTransposeB_CP_4866_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (5) 
      -- CP-element group 59: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_req
      -- CP-element group 59: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/SplitProtocol/$exit
      -- CP-element group 59: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/$exit
      -- CP-element group 59: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/$exit
      -- CP-element group 59: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1797/$exit
      -- 
    phi_stmt_1794_req_5783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1794_req_5783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(59), ack => phi_stmt_1794_req_0); -- 
    convTransposeB_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(57) & convTransposeB_CP_4866_elements(58);
      gj_convTransposeB_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	68 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1638/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(56) & convTransposeB_CP_4866_elements(59);
      gj_convTransposeB_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	53 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/Sample/$exit
      -- 
    ra_5803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1806_inst_ack_0, ack => convTransposeB_CP_4866_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	53 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/Update/ca
      -- 
    ca_5808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1806_inst_ack_1, ack => convTransposeB_CP_4866_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	67 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/SplitProtocol/$exit
      -- CP-element group 63: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/type_cast_1806/$exit
      -- CP-element group 63: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_sources/$exit
      -- CP-element group 63: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/phi_stmt_1800_req
      -- CP-element group 63: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1800/$exit
      -- 
    phi_stmt_1800_req_5809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1800_req_5809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(63), ack => phi_stmt_1800_req_1); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(61) & convTransposeB_CP_4866_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	53 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/Sample/ra
      -- CP-element group 64: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/Sample/$exit
      -- 
    ra_5826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1799_inst_ack_0, ack => convTransposeB_CP_4866_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	53 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/Update/ca
      -- CP-element group 65: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/Update/$exit
      -- 
    ca_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1799_inst_ack_1, ack => convTransposeB_CP_4866_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (5) 
      -- CP-element group 66: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/$exit
      -- CP-element group 66: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/$exit
      -- CP-element group 66: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_req
      -- CP-element group 66: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/phi_stmt_1794_sources/type_cast_1799/SplitProtocol/$exit
      -- CP-element group 66: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1794/$exit
      -- 
    phi_stmt_1794_req_5832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1794_req_5832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(66), ack => phi_stmt_1794_req_1); -- 
    convTransposeB_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(64) & convTransposeB_CP_4866_elements(65);
      gj_convTransposeB_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	63 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1638/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(63) & convTransposeB_CP_4866_elements(66);
      gj_convTransposeB_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  merge  fork  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	60 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1638/merge_stmt_1793_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_1638/merge_stmt_1793_PhiReqMerge
      -- 
    convTransposeB_CP_4866_elements(68) <= OrReduce(convTransposeB_CP_4866_elements(60) & convTransposeB_CP_4866_elements(67));
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1638/merge_stmt_1793_PhiAck/phi_stmt_1794_ack
      -- 
    phi_stmt_1794_ack_5837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1794_ack_0, ack => convTransposeB_CP_4866_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1638/merge_stmt_1793_PhiAck/phi_stmt_1800_ack
      -- 
    phi_stmt_1800_ack_5838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1800_ack_0, ack => convTransposeB_CP_4866_elements(70)); -- 
    -- CP-element group 71:  join  transition  place  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (10) 
      -- CP-element group 71: 	 branch_block_stmt_1638/merge_stmt_1793__exit__
      -- CP-element group 71: 	 branch_block_stmt_1638/assign_stmt_1812_to_assign_stmt_1857__entry__
      -- CP-element group 71: 	 branch_block_stmt_1638/assign_stmt_1812_to_assign_stmt_1857__exit__
      -- CP-element group 71: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 71: 	 branch_block_stmt_1638/assign_stmt_1812_to_assign_stmt_1857/$entry
      -- CP-element group 71: 	 branch_block_stmt_1638/assign_stmt_1812_to_assign_stmt_1857/$exit
      -- CP-element group 71: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1860/$entry
      -- CP-element group 71: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_1638/merge_stmt_1793_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(69) & convTransposeB_CP_4866_elements(70);
      gj_convTransposeB_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Sample/$exit
      -- 
    ra_5858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1863_inst_ack_0, ack => convTransposeB_CP_4866_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	48 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Update/ca
      -- CP-element group 73: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/Update/$exit
      -- 
    ca_5863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1863_inst_ack_1, ack => convTransposeB_CP_4866_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_req
      -- CP-element group 74: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1863/$exit
      -- CP-element group 74: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1860/$exit
      -- CP-element group 74: 	 branch_block_stmt_1638/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1860_req_5864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1860_req_5864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(74), ack => phi_stmt_1860_req_0); -- 
    convTransposeB_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4866_elements(72) & convTransposeB_CP_4866_elements(73);
      gj_convTransposeB_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4866_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_req
      -- CP-element group 75: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/type_cast_1866_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1860/phi_stmt_1860_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1860/$exit
      -- CP-element group 75: 	 branch_block_stmt_1638/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1860_req_5875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1860_req_5875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(75), ack => phi_stmt_1860_req_1); -- 
    -- Element group convTransposeB_CP_4866_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeB_CP_4866_elements(71), ack => convTransposeB_CP_4866_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  merge  transition  place  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1638/merge_stmt_1859_PhiAck/$entry
      -- CP-element group 76: 	 branch_block_stmt_1638/merge_stmt_1859_PhiReqMerge
      -- 
    convTransposeB_CP_4866_elements(76) <= OrReduce(convTransposeB_CP_4866_elements(74) & convTransposeB_CP_4866_elements(75));
    -- CP-element group 77:  fork  transition  place  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	28 
    -- CP-element group 77: 	29 
    -- CP-element group 77: 	31 
    -- CP-element group 77: 	33 
    -- CP-element group 77: 	36 
    -- CP-element group 77: 	37 
    -- CP-element group 77: 	39 
    -- CP-element group 77: 	41 
    -- CP-element group 77: 	44 
    -- CP-element group 77: 	45 
    -- CP-element group 77: 	46 
    -- CP-element group 77: 	35 
    -- CP-element group 77:  members (45) 
      -- CP-element group 77: 	 branch_block_stmt_1638/merge_stmt_1859_PhiAck/$exit
      -- CP-element group 77: 	 branch_block_stmt_1638/merge_stmt_1859_PhiAck/phi_stmt_1860_ack
      -- CP-element group 77: 	 branch_block_stmt_1638/merge_stmt_1859__exit__
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940__entry__
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1886_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_update_start
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1898_final_index_sum_regn_Update/req
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1899_complete/req
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1903_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1907_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_update_start
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/array_obj_ref_1919_final_index_sum_regn_Update/req
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/addr_of_1920_complete/req
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/ptr_deref_1923_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1638/assign_stmt_1873_to_assign_stmt_1940/type_cast_1928_Update/cr
      -- 
    phi_stmt_1860_ack_5880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1860_ack_0, ack => convTransposeB_CP_4866_elements(77)); -- 
    rr_5448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => type_cast_1886_inst_req_0); -- 
    cr_5453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => type_cast_1886_inst_req_1); -- 
    req_5484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => array_obj_ref_1898_index_offset_req_1); -- 
    req_5499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => addr_of_1899_final_reg_req_1); -- 
    cr_5544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => ptr_deref_1903_load_0_req_1); -- 
    rr_5558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => type_cast_1907_inst_req_0); -- 
    cr_5563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => type_cast_1907_inst_req_1); -- 
    req_5594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => array_obj_ref_1919_index_offset_req_1); -- 
    req_5609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => addr_of_1920_final_reg_req_1); -- 
    cr_5659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => ptr_deref_1923_store_0_req_1); -- 
    rr_5668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => type_cast_1928_inst_req_0); -- 
    cr_5673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4866_elements(77), ack => type_cast_1928_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_padding_1696_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1696_word_address_0 : std_logic_vector(0 downto 0);
    signal R_shr114_1897_resized : std_logic_vector(13 downto 0);
    signal R_shr114_1897_scaled : std_logic_vector(13 downto 0);
    signal R_shr67116_1918_resized : std_logic_vector(13 downto 0);
    signal R_shr67116_1918_scaled : std_logic_vector(13 downto 0);
    signal add20_1878 : std_logic_vector(15 downto 0);
    signal add60_1883 : std_logic_vector(15 downto 0);
    signal add73_1935 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1898_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1898_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1898_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1898_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1898_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1898_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1919_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1919_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1919_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1919_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1919_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1919_root_address : std_logic_vector(13 downto 0);
    signal arrayidx69_1921 : std_logic_vector(31 downto 0);
    signal arrayidx_1900 : std_logic_vector(31 downto 0);
    signal call_1641 : std_logic_vector(15 downto 0);
    signal cmp100_1999 : std_logic_vector(0 downto 0);
    signal cmp86_1966 : std_logic_vector(0 downto 0);
    signal cmp_1940 : std_logic_vector(0 downto 0);
    signal conv63_1887 : std_logic_vector(63 downto 0);
    signal conv66_1908 : std_logic_vector(63 downto 0);
    signal conv72_1929 : std_logic_vector(31 downto 0);
    signal conv75_1747 : std_logic_vector(31 downto 0);
    signal conv96_1994 : std_logic_vector(31 downto 0);
    signal conv98_1763 : std_logic_vector(31 downto 0);
    signal div93_1978 : std_logic_vector(15 downto 0);
    signal div99_1769 : std_logic_vector(31 downto 0);
    signal div_1660 : std_logic_vector(15 downto 0);
    signal iNsTr_10_1755 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1650 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1668 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1678 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1690 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1703 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1715 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1727 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1739 : std_logic_vector(31 downto 0);
    signal inc90_1972 : std_logic_vector(15 downto 0);
    signal inc_1961 : std_logic_vector(15 downto 0);
    signal indvar_1860 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1953 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_1990 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1800 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1794 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1984 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1873 : std_logic_vector(15 downto 0);
    signal ptr_deref_1653_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1653_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1653_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1653_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1653_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1671_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1671_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1671_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1671_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1671_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1681_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1681_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1681_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1681_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1681_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1693_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1693_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1693_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1693_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1693_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1706_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1706_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1706_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1706_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1706_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1718_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1718_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1718_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1718_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1718_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1730_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1730_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1730_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1730_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1730_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1742_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1742_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1742_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1742_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1742_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1758_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1758_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1758_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1758_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1758_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1903_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1903_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1903_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1903_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1903_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1923_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1923_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1923_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1923_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1923_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1923_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr114_1893 : std_logic_vector(63 downto 0);
    signal shr67116_1914 : std_logic_vector(63 downto 0);
    signal tmp10_1842 : std_logic_vector(15 downto 0);
    signal tmp11_1672 : std_logic_vector(15 downto 0);
    signal tmp12_1847 : std_logic_vector(15 downto 0);
    signal tmp130_1812 : std_logic_vector(15 downto 0);
    signal tmp131_1817 : std_logic_vector(15 downto 0);
    signal tmp132_1822 : std_logic_vector(15 downto 0);
    signal tmp13_1852 : std_logic_vector(15 downto 0);
    signal tmp14_1857 : std_logic_vector(15 downto 0);
    signal tmp24_1682 : std_logic_vector(15 downto 0);
    signal tmp27_1694 : std_logic_vector(15 downto 0);
    signal tmp30_1697 : std_logic_vector(15 downto 0);
    signal tmp36_1707 : std_logic_vector(15 downto 0);
    signal tmp39_1719 : std_logic_vector(15 downto 0);
    signal tmp3_1775 : std_logic_vector(15 downto 0);
    signal tmp49_1731 : std_logic_vector(15 downto 0);
    signal tmp4_1780 : std_logic_vector(15 downto 0);
    signal tmp53_1743 : std_logic_vector(15 downto 0);
    signal tmp5_1827 : std_logic_vector(15 downto 0);
    signal tmp64_1904 : std_logic_vector(63 downto 0);
    signal tmp6_1832 : std_logic_vector(15 downto 0);
    signal tmp7_1786 : std_logic_vector(15 downto 0);
    signal tmp8_1791 : std_logic_vector(15 downto 0);
    signal tmp97_1759 : std_logic_vector(15 downto 0);
    signal tmp9_1837 : std_logic_vector(15 downto 0);
    signal tmp_1654 : std_logic_vector(15 downto 0);
    signal type_cast_1658_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1767_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1773_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1784_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1797_wire : std_logic_vector(15 downto 0);
    signal type_cast_1799_wire : std_logic_vector(15 downto 0);
    signal type_cast_1804_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1806_wire : std_logic_vector(15 downto 0);
    signal type_cast_1863_wire : std_logic_vector(15 downto 0);
    signal type_cast_1866_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1871_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1891_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1912_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1933_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1951_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1959_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1970_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1976_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_padding_1696_word_address_0 <= "0";
    array_obj_ref_1898_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1898_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1898_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1898_resized_base_address <= "00000000000000";
    array_obj_ref_1919_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1919_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1919_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1919_resized_base_address <= "00000000000000";
    iNsTr_10_1755 <= "00000000000000000000000000000011";
    iNsTr_2_1650 <= "00000000000000000000000000000100";
    iNsTr_3_1668 <= "00000000000000000000000000000101";
    iNsTr_4_1678 <= "00000000000000000000000000000000";
    iNsTr_5_1690 <= "00000000000000000000000000000100";
    iNsTr_6_1703 <= "00000000000000000000000000000001";
    iNsTr_7_1715 <= "00000000000000000000000000000101";
    iNsTr_8_1727 <= "00000000000000000000000000000101";
    iNsTr_9_1739 <= "00000000000000000000000000000100";
    ptr_deref_1653_word_offset_0 <= "0000000";
    ptr_deref_1671_word_offset_0 <= "0000000";
    ptr_deref_1681_word_offset_0 <= "0";
    ptr_deref_1693_word_offset_0 <= "0000000";
    ptr_deref_1706_word_offset_0 <= "0";
    ptr_deref_1718_word_offset_0 <= "0000000";
    ptr_deref_1730_word_offset_0 <= "0000000";
    ptr_deref_1742_word_offset_0 <= "0000000";
    ptr_deref_1758_word_offset_0 <= "0000000";
    ptr_deref_1903_word_offset_0 <= "00000000000000";
    ptr_deref_1923_word_offset_0 <= "00000000000000";
    type_cast_1658_wire_constant <= "0000000000000001";
    type_cast_1767_wire_constant <= "00000000000000000000000000000001";
    type_cast_1773_wire_constant <= "1111111111111111";
    type_cast_1784_wire_constant <= "1111111111111111";
    type_cast_1804_wire_constant <= "0000000000000000";
    type_cast_1866_wire_constant <= "0000000000000000";
    type_cast_1871_wire_constant <= "0000000000000100";
    type_cast_1891_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1912_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1933_wire_constant <= "00000000000000000000000000000100";
    type_cast_1951_wire_constant <= "0000000000000001";
    type_cast_1959_wire_constant <= "0000000000000001";
    type_cast_1970_wire_constant <= "0000000000000001";
    type_cast_1976_wire_constant <= "0000000000000001";
    phi_stmt_1794: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1797_wire & type_cast_1799_wire;
      req <= phi_stmt_1794_req_0 & phi_stmt_1794_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1794",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1794_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1794,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1794
    phi_stmt_1800: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1804_wire_constant & type_cast_1806_wire;
      req <= phi_stmt_1800_req_0 & phi_stmt_1800_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1800",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1800_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1800,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1800
    phi_stmt_1860: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1863_wire & type_cast_1866_wire_constant;
      req <= phi_stmt_1860_req_0 & phi_stmt_1860_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1860",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1860_ack_0,
          idata => idata,
          odata => indvar_1860,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1860
    -- flow-through select operator MUX_1983_inst
    input_dim1x_x2_1984 <= div93_1978 when (cmp86_1966(0) /=  '0') else inc_1961;
    -- flow-through select operator MUX_1989_inst
    input_dim0x_x0_1990 <= inc90_1972 when (cmp86_1966(0) /=  '0') else input_dim0x_x2x_xph_1800;
    addr_of_1899_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1899_final_reg_req_0;
      addr_of_1899_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1899_final_reg_req_1;
      addr_of_1899_final_reg_ack_1<= rack(0);
      addr_of_1899_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1899_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1898_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1900,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1920_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1920_final_reg_req_0;
      addr_of_1920_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1920_final_reg_req_1;
      addr_of_1920_final_reg_ack_1<= rack(0);
      addr_of_1920_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1920_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1919_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx69_1921,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1746_inst_req_0;
      type_cast_1746_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1746_inst_req_1;
      type_cast_1746_inst_ack_1<= rack(0);
      type_cast_1746_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1746_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp11_1672,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_1747,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1762_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1762_inst_req_0;
      type_cast_1762_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1762_inst_req_1;
      type_cast_1762_inst_ack_1<= rack(0);
      type_cast_1762_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1762_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp97_1759,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_1763,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1797_inst_req_0;
      type_cast_1797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1797_inst_req_1;
      type_cast_1797_inst_ack_1<= rack(0);
      type_cast_1797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1797_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1799_inst_req_0;
      type_cast_1799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1799_inst_req_1;
      type_cast_1799_inst_ack_1<= rack(0);
      type_cast_1799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1799_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1806_inst_req_0;
      type_cast_1806_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1806_inst_req_1;
      type_cast_1806_inst_ack_1<= rack(0);
      type_cast_1806_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1806_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_1990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1806_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1863_inst_req_0;
      type_cast_1863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1863_inst_req_1;
      type_cast_1863_inst_ack_1<= rack(0);
      type_cast_1863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1953,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1863_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1886_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1886_inst_req_0;
      type_cast_1886_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1886_inst_req_1;
      type_cast_1886_inst_ack_1<= rack(0);
      type_cast_1886_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1886_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add20_1878,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_1887,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1907_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1907_inst_req_0;
      type_cast_1907_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1907_inst_req_1;
      type_cast_1907_inst_ack_1<= rack(0);
      type_cast_1907_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1907_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add60_1883,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1908,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1928_inst_req_0;
      type_cast_1928_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1928_inst_req_1;
      type_cast_1928_inst_ack_1<= rack(0);
      type_cast_1928_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1873,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_1929,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1993_inst_req_0;
      type_cast_1993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1993_inst_req_1;
      type_cast_1993_inst_ack_1<= rack(0);
      type_cast_1993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_1990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_1994,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1696_gather_scatter
    process(LOAD_padding_1696_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1696_data_0;
      ov(15 downto 0) := iv;
      tmp30_1697 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1898_index_1_rename
    process(R_shr114_1897_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr114_1897_resized;
      ov(13 downto 0) := iv;
      R_shr114_1897_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1898_index_1_resize
    process(shr114_1893) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr114_1893;
      ov := iv(13 downto 0);
      R_shr114_1897_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1898_root_address_inst
    process(array_obj_ref_1898_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1898_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1898_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1919_index_1_rename
    process(R_shr67116_1918_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr67116_1918_resized;
      ov(13 downto 0) := iv;
      R_shr67116_1918_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1919_index_1_resize
    process(shr67116_1914) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr67116_1914;
      ov := iv(13 downto 0);
      R_shr67116_1918_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1919_root_address_inst
    process(array_obj_ref_1919_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1919_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1919_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1653_addr_0
    process(ptr_deref_1653_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1653_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1653_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1653_base_resize
    process(iNsTr_2_1650) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1650;
      ov := iv(6 downto 0);
      ptr_deref_1653_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1653_gather_scatter
    process(ptr_deref_1653_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1653_data_0;
      ov(15 downto 0) := iv;
      tmp_1654 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1653_root_address_inst
    process(ptr_deref_1653_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1653_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1653_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1671_addr_0
    process(ptr_deref_1671_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1671_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1671_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1671_base_resize
    process(iNsTr_3_1668) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1668;
      ov := iv(6 downto 0);
      ptr_deref_1671_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1671_gather_scatter
    process(ptr_deref_1671_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1671_data_0;
      ov(15 downto 0) := iv;
      tmp11_1672 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1671_root_address_inst
    process(ptr_deref_1671_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1671_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1671_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1681_addr_0
    process(ptr_deref_1681_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1681_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1681_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1681_base_resize
    process(iNsTr_4_1678) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1678;
      ov := iv(0 downto 0);
      ptr_deref_1681_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1681_gather_scatter
    process(ptr_deref_1681_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1681_data_0;
      ov(15 downto 0) := iv;
      tmp24_1682 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1681_root_address_inst
    process(ptr_deref_1681_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1681_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1681_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1693_addr_0
    process(ptr_deref_1693_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1693_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1693_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1693_base_resize
    process(iNsTr_5_1690) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1690;
      ov := iv(6 downto 0);
      ptr_deref_1693_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1693_gather_scatter
    process(ptr_deref_1693_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1693_data_0;
      ov(15 downto 0) := iv;
      tmp27_1694 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1693_root_address_inst
    process(ptr_deref_1693_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1693_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1693_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1706_addr_0
    process(ptr_deref_1706_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1706_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1706_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1706_base_resize
    process(iNsTr_6_1703) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1703;
      ov := iv(0 downto 0);
      ptr_deref_1706_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1706_gather_scatter
    process(ptr_deref_1706_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1706_data_0;
      ov(15 downto 0) := iv;
      tmp36_1707 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1706_root_address_inst
    process(ptr_deref_1706_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1706_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1706_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1718_addr_0
    process(ptr_deref_1718_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1718_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1718_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1718_base_resize
    process(iNsTr_7_1715) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1715;
      ov := iv(6 downto 0);
      ptr_deref_1718_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1718_gather_scatter
    process(ptr_deref_1718_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1718_data_0;
      ov(15 downto 0) := iv;
      tmp39_1719 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1718_root_address_inst
    process(ptr_deref_1718_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1718_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1718_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1730_addr_0
    process(ptr_deref_1730_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1730_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1730_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1730_base_resize
    process(iNsTr_8_1727) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1727;
      ov := iv(6 downto 0);
      ptr_deref_1730_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1730_gather_scatter
    process(ptr_deref_1730_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1730_data_0;
      ov(15 downto 0) := iv;
      tmp49_1731 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1730_root_address_inst
    process(ptr_deref_1730_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1730_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1730_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1742_addr_0
    process(ptr_deref_1742_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1742_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1742_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1742_base_resize
    process(iNsTr_9_1739) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1739;
      ov := iv(6 downto 0);
      ptr_deref_1742_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1742_gather_scatter
    process(ptr_deref_1742_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1742_data_0;
      ov(15 downto 0) := iv;
      tmp53_1743 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1742_root_address_inst
    process(ptr_deref_1742_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1742_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1742_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1758_addr_0
    process(ptr_deref_1758_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1758_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1758_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1758_base_resize
    process(iNsTr_10_1755) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1755;
      ov := iv(6 downto 0);
      ptr_deref_1758_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1758_gather_scatter
    process(ptr_deref_1758_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1758_data_0;
      ov(15 downto 0) := iv;
      tmp97_1759 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1758_root_address_inst
    process(ptr_deref_1758_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1758_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1758_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1903_addr_0
    process(ptr_deref_1903_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1903_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1903_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1903_base_resize
    process(arrayidx_1900) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1900;
      ov := iv(13 downto 0);
      ptr_deref_1903_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1903_gather_scatter
    process(ptr_deref_1903_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1903_data_0;
      ov(63 downto 0) := iv;
      tmp64_1904 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1903_root_address_inst
    process(ptr_deref_1903_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1903_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1903_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1923_addr_0
    process(ptr_deref_1923_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1923_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1923_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1923_base_resize
    process(arrayidx69_1921) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx69_1921;
      ov := iv(13 downto 0);
      ptr_deref_1923_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1923_gather_scatter
    process(tmp64_1904) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp64_1904;
      ov(63 downto 0) := iv;
      ptr_deref_1923_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1923_root_address_inst
    process(ptr_deref_1923_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1923_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1923_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1941_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1940;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1941_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1941_branch_req_0,
          ack0 => if_stmt_1941_branch_ack_0,
          ack1 => if_stmt_1941_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2000_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp100_1999;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2000_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2000_branch_req_0,
          ack0 => if_stmt_2000_branch_ack_0,
          ack1 => if_stmt_2000_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1774_inst
    process(tmp39_1719) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp39_1719, type_cast_1773_wire_constant, tmp_var);
      tmp3_1775 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1785_inst
    process(tmp27_1694) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp27_1694, type_cast_1784_wire_constant, tmp_var);
      tmp7_1786 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1816_inst
    process(input_dim1x_x1x_xph_1794, tmp130_1812) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1794, tmp130_1812, tmp_var);
      tmp131_1817 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1831_inst
    process(tmp4_1780, tmp5_1827) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_1780, tmp5_1827, tmp_var);
      tmp6_1832 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1841_inst
    process(tmp8_1791, tmp9_1837) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp8_1791, tmp9_1837, tmp_var);
      tmp10_1842 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1851_inst
    process(tmp6_1832, tmp12_1847) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp6_1832, tmp12_1847, tmp_var);
      tmp13_1852 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1877_inst
    process(tmp132_1822, input_dim2x_x1_1873) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp132_1822, input_dim2x_x1_1873, tmp_var);
      add20_1878 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1882_inst
    process(tmp14_1857, input_dim2x_x1_1873) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_1857, input_dim2x_x1_1873, tmp_var);
      add60_1883 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1952_inst
    process(indvar_1860) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1860, type_cast_1951_wire_constant, tmp_var);
      indvarx_xnext_1953 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1960_inst
    process(input_dim1x_x1x_xph_1794) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1794, type_cast_1959_wire_constant, tmp_var);
      inc_1961 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1971_inst
    process(input_dim0x_x2x_xph_1800) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_1800, type_cast_1970_wire_constant, tmp_var);
      inc90_1972 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1934_inst
    process(conv72_1929) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv72_1929, type_cast_1933_wire_constant, tmp_var);
      add73_1935 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1965_inst
    process(inc_1961, tmp_1654) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1961, tmp_1654, tmp_var);
      cmp86_1966 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1998_inst
    process(conv96_1994, div99_1769) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv96_1994, div99_1769, tmp_var);
      cmp100_1999 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1659_inst
    process(tmp_1654) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1654, type_cast_1658_wire_constant, tmp_var);
      div_1660 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1977_inst
    process(tmp_1654) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1654, type_cast_1976_wire_constant, tmp_var);
      div93_1978 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1768_inst
    process(conv98_1763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv98_1763, type_cast_1767_wire_constant, tmp_var);
      div99_1769 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1892_inst
    process(conv63_1887) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv63_1887, type_cast_1891_wire_constant, tmp_var);
      shr114_1893 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1913_inst
    process(conv66_1908) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv66_1908, type_cast_1912_wire_constant, tmp_var);
      shr67116_1914 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1811_inst
    process(tmp_1654, input_dim0x_x2x_xph_1800) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1654, input_dim0x_x2x_xph_1800, tmp_var);
      tmp130_1812 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1821_inst
    process(tmp11_1672, tmp131_1817) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp11_1672, tmp131_1817, tmp_var);
      tmp132_1822 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1826_inst
    process(tmp36_1707, input_dim1x_x1x_xph_1794) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp36_1707, input_dim1x_x1x_xph_1794, tmp_var);
      tmp5_1827 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1836_inst
    process(tmp24_1682, input_dim0x_x2x_xph_1800) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp24_1682, input_dim0x_x2x_xph_1800, tmp_var);
      tmp9_1837 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1846_inst
    process(tmp53_1743, tmp10_1842) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp53_1743, tmp10_1842, tmp_var);
      tmp12_1847 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1856_inst
    process(tmp49_1731, tmp13_1852) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp49_1731, tmp13_1852, tmp_var);
      tmp14_1857 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1872_inst
    process(indvar_1860) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1860, type_cast_1871_wire_constant, tmp_var);
      input_dim2x_x1_1873 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1779_inst
    process(tmp3_1775, tmp30_1697) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp3_1775, tmp30_1697, tmp_var);
      tmp4_1780 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1790_inst
    process(tmp7_1786, tmp30_1697) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp7_1786, tmp30_1697, tmp_var);
      tmp8_1791 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1939_inst
    process(add73_1935, conv75_1747) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add73_1935, conv75_1747, tmp_var);
      cmp_1940 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_1898_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr114_1897_scaled;
      array_obj_ref_1898_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1898_index_offset_req_0;
      array_obj_ref_1898_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1898_index_offset_req_1;
      array_obj_ref_1898_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_1919_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr67116_1918_scaled;
      array_obj_ref_1919_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1919_index_offset_req_0;
      array_obj_ref_1919_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1919_index_offset_req_1;
      array_obj_ref_1919_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : LOAD_padding_1696_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1696_load_0_req_0;
      LOAD_padding_1696_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1696_load_0_req_1;
      LOAD_padding_1696_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1696_word_address_0;
      LOAD_padding_1696_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1758_load_0 ptr_deref_1653_load_0 ptr_deref_1671_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1758_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1653_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1671_load_0_req_0;
      ptr_deref_1758_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1653_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1671_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1758_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1653_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1671_load_0_req_1;
      ptr_deref_1758_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1653_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1671_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1758_word_address_0 & ptr_deref_1653_word_address_0 & ptr_deref_1671_word_address_0;
      ptr_deref_1758_data_0 <= data_out(47 downto 32);
      ptr_deref_1653_data_0 <= data_out(31 downto 16);
      ptr_deref_1671_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1706_load_0 ptr_deref_1681_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1706_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1681_load_0_req_0;
      ptr_deref_1706_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1681_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1706_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1681_load_0_req_1;
      ptr_deref_1706_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1681_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1706_word_address_0 & ptr_deref_1681_word_address_0;
      ptr_deref_1706_data_0 <= data_out(31 downto 16);
      ptr_deref_1681_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1718_load_0 ptr_deref_1693_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1718_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1693_load_0_req_0;
      ptr_deref_1718_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1693_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1718_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1693_load_0_req_1;
      ptr_deref_1718_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1693_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1718_word_address_0 & ptr_deref_1693_word_address_0;
      ptr_deref_1718_data_0 <= data_out(31 downto 16);
      ptr_deref_1693_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1742_load_0 ptr_deref_1730_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1742_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1730_load_0_req_0;
      ptr_deref_1742_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1730_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1742_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1730_load_0_req_1;
      ptr_deref_1742_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1730_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1742_word_address_0 & ptr_deref_1730_word_address_0;
      ptr_deref_1742_data_0 <= data_out(31 downto 16);
      ptr_deref_1730_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1903_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1903_load_0_req_0;
      ptr_deref_1903_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1903_load_0_req_1;
      ptr_deref_1903_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1903_word_address_0;
      ptr_deref_1903_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1923_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1923_store_0_req_0;
      ptr_deref_1923_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1923_store_0_req_1;
      ptr_deref_1923_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1923_word_address_0;
      data_in <= ptr_deref_1923_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1640_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_start_1640_inst_req_0;
      RPIPE_Block1_start_1640_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_start_1640_inst_req_1;
      RPIPE_Block1_start_1640_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1641 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2008_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2008_inst_req_0;
      WPIPE_Block1_done_2008_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2008_inst_req_1;
      WPIPE_Block1_done_2008_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1641;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5921_start: Boolean;
  signal convTransposeC_CP_5921_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2049_load_0_ack_0 : boolean;
  signal ptr_deref_2071_load_0_req_0 : boolean;
  signal ptr_deref_2049_load_0_req_0 : boolean;
  signal ptr_deref_2031_load_0_ack_1 : boolean;
  signal ptr_deref_2031_load_0_req_0 : boolean;
  signal ptr_deref_2061_load_0_req_0 : boolean;
  signal ptr_deref_2061_load_0_ack_0 : boolean;
  signal ptr_deref_2031_load_0_req_1 : boolean;
  signal ptr_deref_2049_load_0_req_1 : boolean;
  signal ptr_deref_2049_load_0_ack_1 : boolean;
  signal ptr_deref_2071_load_0_ack_0 : boolean;
  signal ptr_deref_2061_load_0_req_1 : boolean;
  signal ptr_deref_2061_load_0_ack_1 : boolean;
  signal ptr_deref_2031_load_0_ack_0 : boolean;
  signal phi_stmt_2238_req_1 : boolean;
  signal type_cast_2184_inst_req_0 : boolean;
  signal type_cast_2184_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2018_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2018_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2018_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2018_inst_ack_1 : boolean;
  signal ptr_deref_2071_load_0_req_1 : boolean;
  signal ptr_deref_2071_load_0_ack_1 : boolean;
  signal ptr_deref_2083_load_0_req_0 : boolean;
  signal ptr_deref_2083_load_0_ack_0 : boolean;
  signal ptr_deref_2083_load_0_req_1 : boolean;
  signal ptr_deref_2083_load_0_ack_1 : boolean;
  signal LOAD_padding_2086_load_0_req_0 : boolean;
  signal LOAD_padding_2086_load_0_ack_0 : boolean;
  signal LOAD_padding_2086_load_0_req_1 : boolean;
  signal LOAD_padding_2086_load_0_ack_1 : boolean;
  signal ptr_deref_2096_load_0_req_0 : boolean;
  signal ptr_deref_2096_load_0_ack_0 : boolean;
  signal ptr_deref_2096_load_0_req_1 : boolean;
  signal ptr_deref_2096_load_0_ack_1 : boolean;
  signal ptr_deref_2108_load_0_req_0 : boolean;
  signal ptr_deref_2108_load_0_ack_0 : boolean;
  signal ptr_deref_2108_load_0_req_1 : boolean;
  signal ptr_deref_2108_load_0_ack_1 : boolean;
  signal ptr_deref_2120_load_0_req_0 : boolean;
  signal ptr_deref_2120_load_0_ack_0 : boolean;
  signal ptr_deref_2120_load_0_req_1 : boolean;
  signal ptr_deref_2120_load_0_ack_1 : boolean;
  signal ptr_deref_2132_load_0_req_0 : boolean;
  signal ptr_deref_2132_load_0_ack_0 : boolean;
  signal ptr_deref_2132_load_0_req_1 : boolean;
  signal ptr_deref_2132_load_0_ack_1 : boolean;
  signal type_cast_2136_inst_req_0 : boolean;
  signal type_cast_2136_inst_ack_0 : boolean;
  signal type_cast_2136_inst_req_1 : boolean;
  signal type_cast_2136_inst_ack_1 : boolean;
  signal phi_stmt_2179_ack_0 : boolean;
  signal type_cast_2140_inst_req_0 : boolean;
  signal type_cast_2140_inst_ack_0 : boolean;
  signal type_cast_2140_inst_req_1 : boolean;
  signal type_cast_2140_inst_ack_1 : boolean;
  signal phi_stmt_2172_ack_0 : boolean;
  signal type_cast_2264_inst_req_0 : boolean;
  signal type_cast_2264_inst_ack_0 : boolean;
  signal type_cast_2264_inst_req_1 : boolean;
  signal type_cast_2264_inst_ack_1 : boolean;
  signal array_obj_ref_2276_index_offset_req_0 : boolean;
  signal array_obj_ref_2276_index_offset_ack_0 : boolean;
  signal array_obj_ref_2276_index_offset_req_1 : boolean;
  signal array_obj_ref_2276_index_offset_ack_1 : boolean;
  signal addr_of_2277_final_reg_req_0 : boolean;
  signal addr_of_2277_final_reg_ack_0 : boolean;
  signal addr_of_2277_final_reg_req_1 : boolean;
  signal addr_of_2277_final_reg_ack_1 : boolean;
  signal type_cast_2244_inst_ack_1 : boolean;
  signal type_cast_2244_inst_req_1 : boolean;
  signal ptr_deref_2281_load_0_req_0 : boolean;
  signal ptr_deref_2281_load_0_ack_0 : boolean;
  signal phi_stmt_2179_req_1 : boolean;
  signal type_cast_2184_inst_ack_1 : boolean;
  signal ptr_deref_2281_load_0_req_1 : boolean;
  signal ptr_deref_2281_load_0_ack_1 : boolean;
  signal type_cast_2184_inst_req_1 : boolean;
  signal type_cast_2285_inst_req_0 : boolean;
  signal type_cast_2285_inst_ack_0 : boolean;
  signal type_cast_2285_inst_req_1 : boolean;
  signal type_cast_2285_inst_ack_1 : boolean;
  signal phi_stmt_2238_ack_0 : boolean;
  signal phi_stmt_2238_req_0 : boolean;
  signal array_obj_ref_2297_index_offset_req_0 : boolean;
  signal array_obj_ref_2297_index_offset_ack_0 : boolean;
  signal array_obj_ref_2297_index_offset_req_1 : boolean;
  signal array_obj_ref_2297_index_offset_ack_1 : boolean;
  signal addr_of_2298_final_reg_req_0 : boolean;
  signal addr_of_2298_final_reg_ack_0 : boolean;
  signal addr_of_2298_final_reg_req_1 : boolean;
  signal addr_of_2298_final_reg_ack_1 : boolean;
  signal type_cast_2244_inst_ack_0 : boolean;
  signal ptr_deref_2301_store_0_req_0 : boolean;
  signal ptr_deref_2301_store_0_ack_0 : boolean;
  signal type_cast_2244_inst_req_0 : boolean;
  signal ptr_deref_2301_store_0_req_1 : boolean;
  signal ptr_deref_2301_store_0_ack_1 : boolean;
  signal type_cast_2306_inst_req_0 : boolean;
  signal type_cast_2306_inst_ack_0 : boolean;
  signal type_cast_2306_inst_req_1 : boolean;
  signal type_cast_2306_inst_ack_1 : boolean;
  signal if_stmt_2319_branch_req_0 : boolean;
  signal if_stmt_2319_branch_ack_1 : boolean;
  signal if_stmt_2319_branch_ack_0 : boolean;
  signal type_cast_2342_inst_req_0 : boolean;
  signal type_cast_2342_inst_ack_0 : boolean;
  signal type_cast_2342_inst_req_1 : boolean;
  signal type_cast_2342_inst_ack_1 : boolean;
  signal type_cast_2351_inst_req_0 : boolean;
  signal type_cast_2351_inst_ack_0 : boolean;
  signal type_cast_2351_inst_req_1 : boolean;
  signal type_cast_2351_inst_ack_1 : boolean;
  signal if_stmt_2370_branch_req_0 : boolean;
  signal if_stmt_2370_branch_ack_1 : boolean;
  signal if_stmt_2370_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2378_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2378_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2378_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2378_inst_ack_1 : boolean;
  signal phi_stmt_2172_req_1 : boolean;
  signal type_cast_2182_inst_req_0 : boolean;
  signal type_cast_2182_inst_ack_0 : boolean;
  signal type_cast_2182_inst_req_1 : boolean;
  signal type_cast_2182_inst_ack_1 : boolean;
  signal phi_stmt_2179_req_0 : boolean;
  signal type_cast_2175_inst_req_0 : boolean;
  signal type_cast_2175_inst_ack_0 : boolean;
  signal type_cast_2175_inst_req_1 : boolean;
  signal type_cast_2175_inst_ack_1 : boolean;
  signal phi_stmt_2172_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5921_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5921_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5921_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5921_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5921: Block -- control-path 
    signal convTransposeC_CP_5921_elements: BooleanArray(79 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5921_elements(0) <= convTransposeC_CP_5921_start;
    convTransposeC_CP_5921_symbol <= convTransposeC_CP_5921_elements(57);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2016/$entry
      -- CP-element group 0: 	 branch_block_stmt_2016/branch_block_stmt_2016__entry__
      -- CP-element group 0: 	 branch_block_stmt_2016/assign_stmt_2019__entry__
      -- CP-element group 0: 	 branch_block_stmt_2016/assign_stmt_2019/$entry
      -- CP-element group 0: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_Sample/rr
      -- 
    rr_5969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(0), ack => RPIPE_Block2_start_2018_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_Update/cr
      -- 
    ra_5970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2018_inst_ack_0, ack => convTransposeC_CP_5921_elements(1)); -- 
    cr_5974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(1), ack => RPIPE_Block2_start_2018_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (259) 
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2019__exit__
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169__entry__
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2019/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2019/RPIPE_Block2_start_2018_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_Update/cr
      -- 
    ca_5975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2018_inst_ack_1, ack => convTransposeC_CP_5921_elements(2)); -- 
    rr_6161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2071_load_0_req_0); -- 
    rr_6061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2049_load_0_req_0); -- 
    rr_6011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2031_load_0_req_0); -- 
    rr_6111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2061_load_0_req_0); -- 
    cr_6022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2031_load_0_req_1); -- 
    cr_6072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2049_load_0_req_1); -- 
    cr_6122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2061_load_0_req_1); -- 
    cr_6172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2071_load_0_req_1); -- 
    rr_6211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2083_load_0_req_0); -- 
    cr_6222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2083_load_0_req_1); -- 
    rr_6244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => LOAD_padding_2086_load_0_req_0); -- 
    cr_6255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => LOAD_padding_2086_load_0_req_1); -- 
    rr_6294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2096_load_0_req_0); -- 
    cr_6305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2096_load_0_req_1); -- 
    rr_6344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2108_load_0_req_0); -- 
    cr_6355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2108_load_0_req_1); -- 
    rr_6394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2120_load_0_req_0); -- 
    cr_6405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2120_load_0_req_1); -- 
    rr_6444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2132_load_0_req_0); -- 
    cr_6455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => ptr_deref_2132_load_0_req_1); -- 
    cr_6474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => type_cast_2136_inst_req_1); -- 
    cr_6488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(2), ack => type_cast_2140_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_sample_completed_
      -- 
    ra_6012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2031_load_0_ack_0, ack => convTransposeC_CP_5921_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	27 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/ptr_deref_2031_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/ptr_deref_2031_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/ptr_deref_2031_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/ptr_deref_2031_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2031_update_completed_
      -- 
    ca_6023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2031_load_0_ack_1, ack => convTransposeC_CP_5921_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Sample/$exit
      -- 
    ra_6062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2049_load_0_ack_0, ack => convTransposeC_CP_5921_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	23 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/ptr_deref_2049_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/ptr_deref_2049_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/ptr_deref_2049_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/ptr_deref_2049_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2049_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_Sample/rr
      -- 
    ca_6073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2049_load_0_ack_1, ack => convTransposeC_CP_5921_elements(6)); -- 
    rr_6469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(6), ack => type_cast_2136_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Sample/word_access_start/$exit
      -- 
    ra_6112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2061_load_0_ack_0, ack => convTransposeC_CP_5921_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	25 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/ptr_deref_2061_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/ptr_deref_2061_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/ptr_deref_2061_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2061_Update/ptr_deref_2061_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_Sample/rr
      -- 
    ca_6123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2061_load_0_ack_1, ack => convTransposeC_CP_5921_elements(8)); -- 
    rr_6483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(8), ack => type_cast_2140_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Sample/word_access_start/word_0/$exit
      -- 
    ra_6162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2071_load_0_ack_0, ack => convTransposeC_CP_5921_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	27 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/ptr_deref_2071_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/ptr_deref_2071_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/ptr_deref_2071_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2071_Update/ptr_deref_2071_Merge/merge_ack
      -- 
    ca_6173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2071_load_0_ack_1, ack => convTransposeC_CP_5921_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Sample/word_access_start/word_0/ra
      -- 
    ra_6212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2083_load_0_ack_0, ack => convTransposeC_CP_5921_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	27 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/ptr_deref_2083_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/ptr_deref_2083_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/ptr_deref_2083_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2083_Update/ptr_deref_2083_Merge/merge_ack
      -- 
    ca_6223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2083_load_0_ack_1, ack => convTransposeC_CP_5921_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Sample/word_access_start/word_0/ra
      -- 
    ra_6245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2086_load_0_ack_0, ack => convTransposeC_CP_5921_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	27 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/LOAD_padding_2086_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/LOAD_padding_2086_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/LOAD_padding_2086_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/LOAD_padding_2086_Update/LOAD_padding_2086_Merge/merge_ack
      -- 
    ca_6256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2086_load_0_ack_1, ack => convTransposeC_CP_5921_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Sample/word_access_start/word_0/ra
      -- 
    ra_6295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2096_load_0_ack_0, ack => convTransposeC_CP_5921_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	27 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/ptr_deref_2096_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/ptr_deref_2096_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/ptr_deref_2096_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2096_Update/ptr_deref_2096_Merge/merge_ack
      -- 
    ca_6306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2096_load_0_ack_1, ack => convTransposeC_CP_5921_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Sample/word_access_start/word_0/ra
      -- 
    ra_6345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2108_load_0_ack_0, ack => convTransposeC_CP_5921_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	27 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/ptr_deref_2108_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/ptr_deref_2108_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/ptr_deref_2108_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2108_Update/ptr_deref_2108_Merge/merge_ack
      -- 
    ca_6356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2108_load_0_ack_1, ack => convTransposeC_CP_5921_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Sample/word_access_start/word_0/ra
      -- 
    ra_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2120_load_0_ack_0, ack => convTransposeC_CP_5921_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	27 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/ptr_deref_2120_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/ptr_deref_2120_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/ptr_deref_2120_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2120_Update/ptr_deref_2120_Merge/merge_ack
      -- 
    ca_6406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2120_load_0_ack_1, ack => convTransposeC_CP_5921_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Sample/word_access_start/word_0/ra
      -- 
    ra_6445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2132_load_0_ack_0, ack => convTransposeC_CP_5921_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/ptr_deref_2132_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/ptr_deref_2132_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/ptr_deref_2132_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/ptr_deref_2132_Update/ptr_deref_2132_Merge/merge_ack
      -- 
    ca_6456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2132_load_0_ack_1, ack => convTransposeC_CP_5921_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	6 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_Sample/ra
      -- 
    ra_6470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2136_inst_ack_0, ack => convTransposeC_CP_5921_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	27 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2136_Update/ca
      -- 
    ca_6475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2136_inst_ack_1, ack => convTransposeC_CP_5921_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	8 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_Sample/ra
      -- 
    ra_6484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2140_inst_ack_0, ack => convTransposeC_CP_5921_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/type_cast_2140_Update/ca
      -- 
    ca_6489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2140_inst_ack_1, ack => convTransposeC_CP_5921_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  place  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	20 
    -- CP-element group 27: 	16 
    -- CP-element group 27: 	12 
    -- CP-element group 27: 	14 
    -- CP-element group 27: 	10 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	24 
    -- CP-element group 27: 	26 
    -- CP-element group 27: 	18 
    -- CP-element group 27: 	4 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	58 
    -- CP-element group 27: 	59 
    -- CP-element group 27: 	60 
    -- CP-element group 27:  members (14) 
      -- CP-element group 27: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169__exit__
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter
      -- CP-element group 27: 	 branch_block_stmt_2016/assign_stmt_2028_to_assign_stmt_2169/$exit
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/Update/cr
      -- 
    rr_6845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(27), ack => type_cast_2182_inst_req_0); -- 
    cr_6850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(27), ack => type_cast_2182_inst_req_1); -- 
    convTransposeC_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(20) & convTransposeC_CP_5921_elements(16) & convTransposeC_CP_5921_elements(12) & convTransposeC_CP_5921_elements(14) & convTransposeC_CP_5921_elements(10) & convTransposeC_CP_5921_elements(22) & convTransposeC_CP_5921_elements(24) & convTransposeC_CP_5921_elements(26) & convTransposeC_CP_5921_elements(18) & convTransposeC_CP_5921_elements(4);
      gj_convTransposeC_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	79 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_Sample/ra
      -- 
    ra_6504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2264_inst_ack_0, ack => convTransposeC_CP_5921_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	79 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (16) 
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_resized_1
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_scaled_1
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_computed_1
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_resize_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_resize_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_resize_1/index_resize_req
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_resize_1/index_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_scale_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_scale_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_scale_1/scale_rename_req
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_index_scale_1/scale_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_Sample/req
      -- 
    ca_6509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2264_inst_ack_1, ack => convTransposeC_CP_5921_elements(29)); -- 
    req_6534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(29), ack => array_obj_ref_2276_index_offset_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	47 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_sample_complete
      -- CP-element group 30: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_Sample/ack
      -- 
    ack_6535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2276_index_offset_ack_0, ack => convTransposeC_CP_5921_elements(30)); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	79 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (11) 
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_offset_calculated
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_request/$entry
      -- CP-element group 31: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_request/req
      -- 
    ack_6540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2276_index_offset_ack_1, ack => convTransposeC_CP_5921_elements(31)); -- 
    req_6549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(31), ack => addr_of_2277_final_reg_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_request/$exit
      -- CP-element group 32: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_request/ack
      -- 
    ack_6550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2277_final_reg_ack_0, ack => convTransposeC_CP_5921_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	79 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (24) 
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_complete/ack
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_word_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_root_address_calculated
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_address_resized
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_addr_resize/$entry
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_addr_resize/$exit
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_addr_resize/base_resize_req
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_addr_resize/base_resize_ack
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_plus_offset/$entry
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_plus_offset/$exit
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_base_plus_offset/sum_rename_ack
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_word_addrgen/$entry
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_word_addrgen/$exit
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_word_addrgen/root_register_req
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_word_addrgen/root_register_ack
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Sample/word_access_start/$entry
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Sample/word_access_start/word_0/$entry
      -- CP-element group 33: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Sample/word_access_start/word_0/rr
      -- 
    ack_6555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2277_final_reg_ack_1, ack => convTransposeC_CP_5921_elements(33)); -- 
    rr_6588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(33), ack => ptr_deref_2281_load_0_req_0); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Sample/word_access_start/$exit
      -- CP-element group 34: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Sample/word_access_start/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Sample/word_access_start/word_0/ra
      -- 
    ra_6589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2281_load_0_ack_0, ack => convTransposeC_CP_5921_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	79 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	42 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/word_access_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/word_access_complete/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/word_access_complete/word_0/ca
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/ptr_deref_2281_Merge/$entry
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/ptr_deref_2281_Merge/$exit
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/ptr_deref_2281_Merge/merge_req
      -- CP-element group 35: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/ptr_deref_2281_Merge/merge_ack
      -- 
    ca_6600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2281_load_0_ack_1, ack => convTransposeC_CP_5921_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	79 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_Sample/ra
      -- 
    ra_6614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2285_inst_ack_0, ack => convTransposeC_CP_5921_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	79 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_resized_1
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_scaled_1
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_computed_1
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_resize_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_resize_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_resize_1/index_resize_req
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_resize_1/index_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_scale_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_scale_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_scale_1/scale_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_index_scale_1/scale_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_Sample/req
      -- 
    ca_6619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2285_inst_ack_1, ack => convTransposeC_CP_5921_elements(37)); -- 
    req_6644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(37), ack => array_obj_ref_2297_index_offset_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_sample_complete
      -- CP-element group 38: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_Sample/ack
      -- 
    ack_6645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2297_index_offset_ack_0, ack => convTransposeC_CP_5921_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	79 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (11) 
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_offset_calculated
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_request/$entry
      -- CP-element group 39: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_request/req
      -- 
    ack_6650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2297_index_offset_ack_1, ack => convTransposeC_CP_5921_elements(39)); -- 
    req_6659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(39), ack => addr_of_2298_final_reg_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_request/$exit
      -- CP-element group 40: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_request/ack
      -- 
    ack_6660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2298_final_reg_ack_0, ack => convTransposeC_CP_5921_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	79 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (19) 
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_complete/ack
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_word_addrgen/root_register_ack
      -- 
    ack_6665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2298_final_reg_ack_1, ack => convTransposeC_CP_5921_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	35 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/ptr_deref_2301_Split/$entry
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/ptr_deref_2301_Split/$exit
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/ptr_deref_2301_Split/split_req
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/ptr_deref_2301_Split/split_ack
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/word_access_start/word_0/rr
      -- 
    rr_6703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(42), ack => ptr_deref_2301_store_0_req_0); -- 
    convTransposeC_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(41) & convTransposeC_CP_5921_elements(35);
      gj_convTransposeC_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Sample/word_access_start/word_0/ra
      -- 
    ra_6704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2301_store_0_ack_0, ack => convTransposeC_CP_5921_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	79 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Update/word_access_complete/word_0/ca
      -- 
    ca_6715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2301_store_0_ack_1, ack => convTransposeC_CP_5921_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	79 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_Sample/ra
      -- 
    ra_6724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_0, ack => convTransposeC_CP_5921_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	79 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_Update/ca
      -- 
    ca_6729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2306_inst_ack_1, ack => convTransposeC_CP_5921_elements(46)); -- 
    -- CP-element group 47:  branch  join  transition  place  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: 	30 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (10) 
      -- CP-element group 47: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318__exit__
      -- CP-element group 47: 	 branch_block_stmt_2016/if_stmt_2319__entry__
      -- CP-element group 47: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/$exit
      -- CP-element group 47: 	 branch_block_stmt_2016/if_stmt_2319_dead_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_2016/if_stmt_2319_eval_test/$entry
      -- CP-element group 47: 	 branch_block_stmt_2016/if_stmt_2319_eval_test/$exit
      -- CP-element group 47: 	 branch_block_stmt_2016/if_stmt_2319_eval_test/branch_req
      -- CP-element group 47: 	 branch_block_stmt_2016/R_cmp_2320_place
      -- CP-element group 47: 	 branch_block_stmt_2016/if_stmt_2319_if_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_2016/if_stmt_2319_else_link/$entry
      -- 
    branch_req_6737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(47), ack => if_stmt_2319_branch_req_0); -- 
    convTransposeC_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(38) & convTransposeC_CP_5921_elements(44) & convTransposeC_CP_5921_elements(46) & convTransposeC_CP_5921_elements(30);
      gj_convTransposeC_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48: 	75 
    -- CP-element group 48:  members (24) 
      -- CP-element group 48: 	 branch_block_stmt_2016/merge_stmt_2325_PhiReqMerge
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/merge_stmt_2325__exit__
      -- CP-element group 48: 	 branch_block_stmt_2016/assign_stmt_2331__entry__
      -- CP-element group 48: 	 branch_block_stmt_2016/assign_stmt_2331__exit__
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/merge_stmt_2325_PhiAck/dummy
      -- CP-element group 48: 	 branch_block_stmt_2016/merge_stmt_2325_PhiAck/$exit
      -- CP-element group 48: 	 branch_block_stmt_2016/merge_stmt_2325_PhiAck/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/Update/cr
      -- CP-element group 48: 	 branch_block_stmt_2016/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_2016/if_stmt_2319_if_link/$exit
      -- CP-element group 48: 	 branch_block_stmt_2016/if_stmt_2319_if_link/if_choice_transition
      -- CP-element group 48: 	 branch_block_stmt_2016/whilex_xbody_ifx_xthen
      -- CP-element group 48: 	 branch_block_stmt_2016/assign_stmt_2331/$entry
      -- CP-element group 48: 	 branch_block_stmt_2016/assign_stmt_2331/$exit
      -- 
    if_choice_transition_6742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2319_branch_ack_1, ack => convTransposeC_CP_5921_elements(48)); -- 
    cr_6931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(48), ack => type_cast_2244_inst_req_1); -- 
    rr_6926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(48), ack => type_cast_2244_inst_req_0); -- 
    -- CP-element group 49:  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	53 
    -- CP-element group 49:  members (21) 
      -- CP-element group 49: 	 branch_block_stmt_2016/merge_stmt_2333_PhiReqMerge
      -- CP-element group 49: 	 branch_block_stmt_2016/merge_stmt_2333__exit__
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369__entry__
      -- CP-element group 49: 	 branch_block_stmt_2016/merge_stmt_2333_PhiAck/dummy
      -- CP-element group 49: 	 branch_block_stmt_2016/merge_stmt_2333_PhiAck/$exit
      -- CP-element group 49: 	 branch_block_stmt_2016/merge_stmt_2333_PhiAck/$entry
      -- CP-element group 49: 	 branch_block_stmt_2016/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 49: 	 branch_block_stmt_2016/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_2016/if_stmt_2319_else_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_2016/if_stmt_2319_else_link/else_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_2016/whilex_xbody_ifx_xelse
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/$entry
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_update_start_
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_update_start_
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_Update/cr
      -- 
    else_choice_transition_6746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2319_branch_ack_0, ack => convTransposeC_CP_5921_elements(49)); -- 
    rr_6762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(49), ack => type_cast_2342_inst_req_0); -- 
    cr_6767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(49), ack => type_cast_2342_inst_req_1); -- 
    cr_6781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(49), ack => type_cast_2351_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_Sample/ra
      -- 
    ra_6763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2342_inst_ack_0, ack => convTransposeC_CP_5921_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2342_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_Sample/rr
      -- 
    ca_6768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2342_inst_ack_1, ack => convTransposeC_CP_5921_elements(51)); -- 
    rr_6776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(51), ack => type_cast_2351_inst_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_Sample/ra
      -- 
    ra_6777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_0, ack => convTransposeC_CP_5921_elements(52)); -- 
    -- CP-element group 53:  branch  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	49 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (13) 
      -- CP-element group 53: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369__exit__
      -- CP-element group 53: 	 branch_block_stmt_2016/if_stmt_2370__entry__
      -- CP-element group 53: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/$exit
      -- CP-element group 53: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2016/assign_stmt_2339_to_assign_stmt_2369/type_cast_2351_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_2016/if_stmt_2370_dead_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2016/if_stmt_2370_eval_test/$entry
      -- CP-element group 53: 	 branch_block_stmt_2016/if_stmt_2370_eval_test/$exit
      -- CP-element group 53: 	 branch_block_stmt_2016/if_stmt_2370_eval_test/branch_req
      -- CP-element group 53: 	 branch_block_stmt_2016/R_cmp97_2371_place
      -- CP-element group 53: 	 branch_block_stmt_2016/if_stmt_2370_if_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_2016/if_stmt_2370_else_link/$entry
      -- 
    ca_6782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2351_inst_ack_1, ack => convTransposeC_CP_5921_elements(53)); -- 
    branch_req_6790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(53), ack => if_stmt_2370_branch_req_0); -- 
    -- CP-element group 54:  merge  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (15) 
      -- CP-element group 54: 	 branch_block_stmt_2016/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_2016/merge_stmt_2376_PhiReqMerge
      -- CP-element group 54: 	 branch_block_stmt_2016/merge_stmt_2376_PhiAck/$entry
      -- CP-element group 54: 	 branch_block_stmt_2016/merge_stmt_2376_PhiAck/$exit
      -- CP-element group 54: 	 branch_block_stmt_2016/merge_stmt_2376_PhiAck/dummy
      -- CP-element group 54: 	 branch_block_stmt_2016/merge_stmt_2376__exit__
      -- CP-element group 54: 	 branch_block_stmt_2016/assign_stmt_2380__entry__
      -- CP-element group 54: 	 branch_block_stmt_2016/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_2016/if_stmt_2370_if_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_2016/if_stmt_2370_if_link/if_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_2016/ifx_xelse_whilex_xend
      -- CP-element group 54: 	 branch_block_stmt_2016/assign_stmt_2380/$entry
      -- CP-element group 54: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_Sample/req
      -- 
    if_choice_transition_6795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2370_branch_ack_1, ack => convTransposeC_CP_5921_elements(54)); -- 
    req_6812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(54), ack => WPIPE_Block2_done_2378_inst_req_0); -- 
    -- CP-element group 55:  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	63 
    -- CP-element group 55: 	64 
    -- CP-element group 55: 	66 
    -- CP-element group 55: 	67 
    -- CP-element group 55:  members (20) 
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/if_stmt_2370_else_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_2016/if_stmt_2370_else_link/else_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/$entry
      -- 
    else_choice_transition_6799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2370_branch_ack_0, ack => convTransposeC_CP_5921_elements(55)); -- 
    rr_6894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(55), ack => type_cast_2184_inst_req_0); -- 
    cr_6899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(55), ack => type_cast_2184_inst_req_1); -- 
    rr_6871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(55), ack => type_cast_2175_inst_req_0); -- 
    cr_6876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(55), ack => type_cast_2175_inst_req_1); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_update_start_
      -- CP-element group 56: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_Sample/ack
      -- CP-element group 56: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_Update/req
      -- 
    ack_6813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2378_inst_ack_0, ack => convTransposeC_CP_5921_elements(56)); -- 
    req_6817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(56), ack => WPIPE_Block2_done_2378_inst_req_1); -- 
    -- CP-element group 57:  transition  place  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (16) 
      -- CP-element group 57: 	 branch_block_stmt_2016/merge_stmt_2382_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_2016/return___PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_2016/return___PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_2016/merge_stmt_2382_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_2016/merge_stmt_2382_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_2016/merge_stmt_2382_PhiAck/dummy
      -- CP-element group 57: 	 $exit
      -- CP-element group 57: 	 branch_block_stmt_2016/$exit
      -- CP-element group 57: 	 branch_block_stmt_2016/branch_block_stmt_2016__exit__
      -- CP-element group 57: 	 branch_block_stmt_2016/assign_stmt_2380__exit__
      -- CP-element group 57: 	 branch_block_stmt_2016/return__
      -- CP-element group 57: 	 branch_block_stmt_2016/merge_stmt_2382__exit__
      -- CP-element group 57: 	 branch_block_stmt_2016/assign_stmt_2380/$exit
      -- CP-element group 57: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2016/assign_stmt_2380/WPIPE_Block2_done_2378_Update/ack
      -- 
    ack_6818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2378_inst_ack_1, ack => convTransposeC_CP_5921_elements(57)); -- 
    -- CP-element group 58:  transition  output  delay-element  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	27 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	62 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/$exit
      -- CP-element group 58: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/$exit
      -- CP-element group 58: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2178_konst_delay_trans
      -- CP-element group 58: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_req
      -- 
    phi_stmt_2172_req_6829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2172_req_6829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(58), ack => phi_stmt_2172_req_1); -- 
    -- Element group convTransposeC_CP_5921_elements(58) is a control-delay.
    cp_element_58_delay: control_delay_element  generic map(name => " 58_delay", delay_value => 1)  port map(req => convTransposeC_CP_5921_elements(27), ack => convTransposeC_CP_5921_elements(58), clk => clk, reset =>reset);
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	27 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/Sample/ra
      -- 
    ra_6846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2182_inst_ack_0, ack => convTransposeC_CP_5921_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/Update/ca
      -- 
    ca_6851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2182_inst_ack_1, ack => convTransposeC_CP_5921_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/$exit
      -- CP-element group 61: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/$exit
      -- CP-element group 61: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/$exit
      -- CP-element group 61: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2182/SplitProtocol/$exit
      -- CP-element group 61: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_req
      -- 
    phi_stmt_2179_req_6852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2179_req_6852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(61), ack => phi_stmt_2179_req_0); -- 
    convTransposeC_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(59) & convTransposeC_CP_5921_elements(60);
      gj_convTransposeC_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	58 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	70 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_2016/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(58) & convTransposeC_CP_5921_elements(61);
      gj_convTransposeC_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	55 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/Sample/ra
      -- 
    ra_6872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2175_inst_ack_0, ack => convTransposeC_CP_5921_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	55 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/Update/ca
      -- 
    ca_6877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2175_inst_ack_1, ack => convTransposeC_CP_5921_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	69 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/$exit
      -- CP-element group 65: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/$exit
      -- CP-element group 65: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_sources/type_cast_2175/SplitProtocol/$exit
      -- CP-element group 65: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2172/phi_stmt_2172_req
      -- 
    phi_stmt_2172_req_6878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2172_req_6878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(65), ack => phi_stmt_2172_req_0); -- 
    convTransposeC_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(63) & convTransposeC_CP_5921_elements(64);
      gj_convTransposeC_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	55 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/Sample/ra
      -- 
    ra_6895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2184_inst_ack_0, ack => convTransposeC_CP_5921_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	55 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/Update/ca
      -- CP-element group 67: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/Update/$exit
      -- 
    ca_6900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2184_inst_ack_1, ack => convTransposeC_CP_5921_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/$exit
      -- CP-element group 68: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/type_cast_2184/SplitProtocol/$exit
      -- CP-element group 68: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_sources/$exit
      -- CP-element group 68: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/phi_stmt_2179_req
      -- CP-element group 68: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2179/$exit
      -- 
    phi_stmt_2179_req_6901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2179_req_6901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(68), ack => phi_stmt_2179_req_1); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(66) & convTransposeC_CP_5921_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	65 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_2016/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(65) & convTransposeC_CP_5921_elements(68);
      gj_convTransposeC_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  merge  fork  transition  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: 	62 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2016/merge_stmt_2171_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2016/merge_stmt_2171_PhiReqMerge
      -- 
    convTransposeC_CP_5921_elements(70) <= OrReduce(convTransposeC_CP_5921_elements(69) & convTransposeC_CP_5921_elements(62));
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2016/merge_stmt_2171_PhiAck/phi_stmt_2172_ack
      -- 
    phi_stmt_2172_ack_6906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2172_ack_0, ack => convTransposeC_CP_5921_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_2016/merge_stmt_2171_PhiAck/phi_stmt_2179_ack
      -- 
    phi_stmt_2179_ack_6907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2179_ack_0, ack => convTransposeC_CP_5921_elements(72)); -- 
    -- CP-element group 73:  join  transition  place  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (10) 
      -- CP-element group 73: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 73: 	 branch_block_stmt_2016/merge_stmt_2171__exit__
      -- CP-element group 73: 	 branch_block_stmt_2016/assign_stmt_2190_to_assign_stmt_2235__entry__
      -- CP-element group 73: 	 branch_block_stmt_2016/assign_stmt_2190_to_assign_stmt_2235__exit__
      -- CP-element group 73: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 73: 	 branch_block_stmt_2016/merge_stmt_2171_PhiAck/$exit
      -- CP-element group 73: 	 branch_block_stmt_2016/assign_stmt_2190_to_assign_stmt_2235/$entry
      -- CP-element group 73: 	 branch_block_stmt_2016/assign_stmt_2190_to_assign_stmt_2235/$exit
      -- CP-element group 73: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/$entry
      -- CP-element group 73: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2238/$entry
      -- 
    convTransposeC_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(71) & convTransposeC_CP_5921_elements(72);
      gj_convTransposeC_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	48 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/Sample/ra
      -- 
    ra_6927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2244_inst_ack_0, ack => convTransposeC_CP_5921_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	48 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/Update/ca
      -- CP-element group 75: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/Update/$exit
      -- 
    ca_6932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2244_inst_ack_1, ack => convTransposeC_CP_5921_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 76: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/$exit
      -- CP-element group 76: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_req
      -- CP-element group 76: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2244/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2016/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2238/$exit
      -- 
    phi_stmt_2238_req_6933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2238_req_6933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(76), ack => phi_stmt_2238_req_1); -- 
    convTransposeC_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5921_elements(74) & convTransposeC_CP_5921_elements(75);
      gj_convTransposeC_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5921_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_req
      -- CP-element group 77: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2238/phi_stmt_2238_sources/type_cast_2242_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2238/$exit
      -- CP-element group 77: 	 branch_block_stmt_2016/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_2238_req_6944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2238_req_6944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(77), ack => phi_stmt_2238_req_0); -- 
    -- Element group convTransposeC_CP_5921_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeC_CP_5921_elements(73), ack => convTransposeC_CP_5921_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  merge  transition  place  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2016/merge_stmt_2237_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2016/merge_stmt_2237_PhiAck/$entry
      -- 
    convTransposeC_CP_5921_elements(78) <= OrReduce(convTransposeC_CP_5921_elements(76) & convTransposeC_CP_5921_elements(77));
    -- CP-element group 79:  fork  transition  place  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	39 
    -- CP-element group 79: 	44 
    -- CP-element group 79: 	45 
    -- CP-element group 79: 	41 
    -- CP-element group 79: 	35 
    -- CP-element group 79: 	46 
    -- CP-element group 79: 	36 
    -- CP-element group 79: 	37 
    -- CP-element group 79: 	28 
    -- CP-element group 79: 	29 
    -- CP-element group 79: 	31 
    -- CP-element group 79: 	33 
    -- CP-element group 79:  members (45) 
      -- CP-element group 79: 	 branch_block_stmt_2016/merge_stmt_2237__exit__
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318__entry__
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2264_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_update_start
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2276_final_index_sum_regn_Update/req
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2277_complete/req
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/word_access_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/word_access_complete/word_0/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2281_Update/word_access_complete/word_0/cr
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2285_Update/cr
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/merge_stmt_2237_PhiAck/phi_stmt_2238_ack
      -- CP-element group 79: 	 branch_block_stmt_2016/merge_stmt_2237_PhiAck/$exit
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_update_start
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/array_obj_ref_2297_final_index_sum_regn_Update/req
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/addr_of_2298_complete/req
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Update/word_access_complete/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Update/word_access_complete/word_0/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/ptr_deref_2301_Update/word_access_complete/word_0/cr
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2016/assign_stmt_2251_to_assign_stmt_2318/type_cast_2306_Update/cr
      -- 
    phi_stmt_2238_ack_6949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2238_ack_0, ack => convTransposeC_CP_5921_elements(79)); -- 
    rr_6503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => type_cast_2264_inst_req_0); -- 
    cr_6508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => type_cast_2264_inst_req_1); -- 
    req_6539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => array_obj_ref_2276_index_offset_req_1); -- 
    req_6554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => addr_of_2277_final_reg_req_1); -- 
    cr_6599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => ptr_deref_2281_load_0_req_1); -- 
    rr_6613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => type_cast_2285_inst_req_0); -- 
    cr_6618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => type_cast_2285_inst_req_1); -- 
    req_6649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => array_obj_ref_2297_index_offset_req_1); -- 
    req_6664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => addr_of_2298_final_reg_req_1); -- 
    cr_6714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => ptr_deref_2301_store_0_req_1); -- 
    rr_6723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => type_cast_2306_inst_req_0); -- 
    cr_6728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5921_elements(79), ack => type_cast_2306_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_padding_2086_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2086_word_address_0 : std_logic_vector(0 downto 0);
    signal R_shr111_2275_resized : std_logic_vector(13 downto 0);
    signal R_shr111_2275_scaled : std_logic_vector(13 downto 0);
    signal R_shr68113_2296_resized : std_logic_vector(13 downto 0);
    signal R_shr68113_2296_scaled : std_logic_vector(13 downto 0);
    signal add21_2256 : std_logic_vector(15 downto 0);
    signal add61_2261 : std_logic_vector(15 downto 0);
    signal add74_2313 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2276_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2276_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2276_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2276_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2276_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2276_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2297_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2297_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2297_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2297_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2297_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2297_root_address : std_logic_vector(13 downto 0);
    signal arrayidx70_2299 : std_logic_vector(31 downto 0);
    signal arrayidx_2278 : std_logic_vector(31 downto 0);
    signal call_2019 : std_logic_vector(15 downto 0);
    signal cmp88_2348 : std_logic_vector(0 downto 0);
    signal cmp97_2369 : std_logic_vector(0 downto 0);
    signal cmp_2318 : std_logic_vector(0 downto 0);
    signal conv64_2265 : std_logic_vector(63 downto 0);
    signal conv67_2286 : std_logic_vector(63 downto 0);
    signal conv73_2307 : std_logic_vector(31 downto 0);
    signal conv76_2137 : std_logic_vector(31 downto 0);
    signal conv84_2343 : std_logic_vector(31 downto 0);
    signal conv86_2141 : std_logic_vector(31 downto 0);
    signal div87_2147 : std_logic_vector(31 downto 0);
    signal div_2038 : std_logic_vector(15 downto 0);
    signal iNsTr_10_2129 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2028 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2046 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2058 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2068 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2080 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2093 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2105 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2117 : std_logic_vector(31 downto 0);
    signal inc92_2352 : std_logic_vector(15 downto 0);
    signal inc92x_xinput_dim0x_x2_2357 : std_logic_vector(15 downto 0);
    signal inc_2339 : std_logic_vector(15 downto 0);
    signal indvar_2238 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2331 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2179 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2172 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2364 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2251 : std_logic_vector(15 downto 0);
    signal ptr_deref_2031_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2031_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2031_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2031_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2031_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2049_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2049_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2049_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2049_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2049_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2061_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2061_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2061_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2061_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2061_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2071_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2071_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2071_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2071_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2071_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2083_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2083_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2083_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2083_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2083_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2096_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2096_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2096_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2096_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2096_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2108_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2108_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2108_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2108_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2108_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2120_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2120_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2120_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2120_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2120_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2132_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2132_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2132_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2132_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2132_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2281_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2281_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2281_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2281_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2281_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2301_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2301_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2301_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2301_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2301_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2301_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr111_2271 : std_logic_vector(63 downto 0);
    signal shr68113_2292 : std_logic_vector(63 downto 0);
    signal tmp10_2220 : std_logic_vector(15 downto 0);
    signal tmp11_2225 : std_logic_vector(15 downto 0);
    signal tmp127_2190 : std_logic_vector(15 downto 0);
    signal tmp128_2195 : std_logic_vector(15 downto 0);
    signal tmp129_2200 : std_logic_vector(15 downto 0);
    signal tmp12_2050 : std_logic_vector(15 downto 0);
    signal tmp13_2230 : std_logic_vector(15 downto 0);
    signal tmp14_2235 : std_logic_vector(15 downto 0);
    signal tmp16_2062 : std_logic_vector(15 downto 0);
    signal tmp25_2072 : std_logic_vector(15 downto 0);
    signal tmp28_2084 : std_logic_vector(15 downto 0);
    signal tmp31_2087 : std_logic_vector(15 downto 0);
    signal tmp37_2097 : std_logic_vector(15 downto 0);
    signal tmp3_2153 : std_logic_vector(15 downto 0);
    signal tmp40_2109 : std_logic_vector(15 downto 0);
    signal tmp4_2158 : std_logic_vector(15 downto 0);
    signal tmp50_2121 : std_logic_vector(15 downto 0);
    signal tmp54_2133 : std_logic_vector(15 downto 0);
    signal tmp5_2205 : std_logic_vector(15 downto 0);
    signal tmp65_2282 : std_logic_vector(63 downto 0);
    signal tmp6_2210 : std_logic_vector(15 downto 0);
    signal tmp7_2164 : std_logic_vector(15 downto 0);
    signal tmp8_2169 : std_logic_vector(15 downto 0);
    signal tmp9_2215 : std_logic_vector(15 downto 0);
    signal tmp_2032 : std_logic_vector(15 downto 0);
    signal type_cast_2036_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2145_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2151_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2162_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2175_wire : std_logic_vector(15 downto 0);
    signal type_cast_2178_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2182_wire : std_logic_vector(15 downto 0);
    signal type_cast_2184_wire : std_logic_vector(15 downto 0);
    signal type_cast_2242_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2244_wire : std_logic_vector(15 downto 0);
    signal type_cast_2249_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2269_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2290_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2311_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2329_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2337_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2361_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_padding_2086_word_address_0 <= "0";
    array_obj_ref_2276_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2276_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2276_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2276_resized_base_address <= "00000000000000";
    array_obj_ref_2297_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2297_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2297_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2297_resized_base_address <= "00000000000000";
    iNsTr_10_2129 <= "00000000000000000000000000000100";
    iNsTr_2_2028 <= "00000000000000000000000000000011";
    iNsTr_3_2046 <= "00000000000000000000000000000101";
    iNsTr_4_2058 <= "00000000000000000000000000000100";
    iNsTr_5_2068 <= "00000000000000000000000000000000";
    iNsTr_6_2080 <= "00000000000000000000000000000100";
    iNsTr_7_2093 <= "00000000000000000000000000000001";
    iNsTr_8_2105 <= "00000000000000000000000000000101";
    iNsTr_9_2117 <= "00000000000000000000000000000101";
    ptr_deref_2031_word_offset_0 <= "0000000";
    ptr_deref_2049_word_offset_0 <= "0000000";
    ptr_deref_2061_word_offset_0 <= "0000000";
    ptr_deref_2071_word_offset_0 <= "0";
    ptr_deref_2083_word_offset_0 <= "0000000";
    ptr_deref_2096_word_offset_0 <= "0";
    ptr_deref_2108_word_offset_0 <= "0000000";
    ptr_deref_2120_word_offset_0 <= "0000000";
    ptr_deref_2132_word_offset_0 <= "0000000";
    ptr_deref_2281_word_offset_0 <= "00000000000000";
    ptr_deref_2301_word_offset_0 <= "00000000000000";
    type_cast_2036_wire_constant <= "0000000000000001";
    type_cast_2145_wire_constant <= "00000000000000000000000000000001";
    type_cast_2151_wire_constant <= "1111111111111111";
    type_cast_2162_wire_constant <= "1111111111111111";
    type_cast_2178_wire_constant <= "0000000000000000";
    type_cast_2242_wire_constant <= "0000000000000000";
    type_cast_2249_wire_constant <= "0000000000000100";
    type_cast_2269_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2290_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2311_wire_constant <= "00000000000000000000000000000100";
    type_cast_2329_wire_constant <= "0000000000000001";
    type_cast_2337_wire_constant <= "0000000000000001";
    type_cast_2361_wire_constant <= "0000000000000000";
    phi_stmt_2172: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2175_wire & type_cast_2178_wire_constant;
      req <= phi_stmt_2172_req_0 & phi_stmt_2172_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2172",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2172_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2172,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2172
    phi_stmt_2179: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2182_wire & type_cast_2184_wire;
      req <= phi_stmt_2179_req_0 & phi_stmt_2179_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2179",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2179_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2179,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2179
    phi_stmt_2238: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2242_wire_constant & type_cast_2244_wire;
      req <= phi_stmt_2238_req_0 & phi_stmt_2238_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2238",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2238_ack_0,
          idata => idata,
          odata => indvar_2238,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2238
    -- flow-through select operator MUX_2363_inst
    input_dim1x_x2_2364 <= type_cast_2361_wire_constant when (cmp88_2348(0) /=  '0') else inc_2339;
    addr_of_2277_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2277_final_reg_req_0;
      addr_of_2277_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2277_final_reg_req_1;
      addr_of_2277_final_reg_ack_1<= rack(0);
      addr_of_2277_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2277_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2276_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2278,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2298_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2298_final_reg_req_0;
      addr_of_2298_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2298_final_reg_req_1;
      addr_of_2298_final_reg_ack_1<= rack(0);
      addr_of_2298_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2298_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2297_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx70_2299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2136_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2136_inst_req_0;
      type_cast_2136_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2136_inst_req_1;
      type_cast_2136_inst_ack_1<= rack(0);
      type_cast_2136_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2136_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_2050,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2137,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2140_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2140_inst_req_0;
      type_cast_2140_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2140_inst_req_1;
      type_cast_2140_inst_ack_1<= rack(0);
      type_cast_2140_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2140_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp16_2062,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2141,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2175_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2175_inst_req_0;
      type_cast_2175_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2175_inst_req_1;
      type_cast_2175_inst_ack_1<= rack(0);
      type_cast_2175_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2175_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2364,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2175_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2182_inst_req_0;
      type_cast_2182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2182_inst_req_1;
      type_cast_2182_inst_ack_1<= rack(0);
      type_cast_2182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2038,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2182_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2184_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2184_inst_req_0;
      type_cast_2184_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2184_inst_req_1;
      type_cast_2184_inst_ack_1<= rack(0);
      type_cast_2184_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2184_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc92x_xinput_dim0x_x2_2357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2184_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2244_inst_req_0;
      type_cast_2244_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2244_inst_req_1;
      type_cast_2244_inst_ack_1<= rack(0);
      type_cast_2244_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2244_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2331,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2244_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2264_inst_req_0;
      type_cast_2264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2264_inst_req_1;
      type_cast_2264_inst_ack_1<= rack(0);
      type_cast_2264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_2256,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_2265,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2285_inst_req_0;
      type_cast_2285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2285_inst_req_1;
      type_cast_2285_inst_ack_1<= rack(0);
      type_cast_2285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add61_2261,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_2286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2306_inst_req_0;
      type_cast_2306_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2306_inst_req_1;
      type_cast_2306_inst_ack_1<= rack(0);
      type_cast_2306_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2307,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2342_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2342_inst_req_0;
      type_cast_2342_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2342_inst_req_1;
      type_cast_2342_inst_ack_1<= rack(0);
      type_cast_2342_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2342_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2343,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2351_inst_req_0;
      type_cast_2351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2351_inst_req_1;
      type_cast_2351_inst_ack_1<= rack(0);
      type_cast_2351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp88_2348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc92_2352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2086_gather_scatter
    process(LOAD_padding_2086_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2086_data_0;
      ov(15 downto 0) := iv;
      tmp31_2087 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2276_index_1_rename
    process(R_shr111_2275_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr111_2275_resized;
      ov(13 downto 0) := iv;
      R_shr111_2275_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2276_index_1_resize
    process(shr111_2271) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr111_2271;
      ov := iv(13 downto 0);
      R_shr111_2275_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2276_root_address_inst
    process(array_obj_ref_2276_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2276_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2276_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2297_index_1_rename
    process(R_shr68113_2296_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr68113_2296_resized;
      ov(13 downto 0) := iv;
      R_shr68113_2296_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2297_index_1_resize
    process(shr68113_2292) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr68113_2292;
      ov := iv(13 downto 0);
      R_shr68113_2296_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2297_root_address_inst
    process(array_obj_ref_2297_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2297_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2297_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2031_addr_0
    process(ptr_deref_2031_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2031_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2031_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2031_base_resize
    process(iNsTr_2_2028) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2028;
      ov := iv(6 downto 0);
      ptr_deref_2031_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2031_gather_scatter
    process(ptr_deref_2031_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2031_data_0;
      ov(15 downto 0) := iv;
      tmp_2032 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2031_root_address_inst
    process(ptr_deref_2031_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2031_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2031_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2049_addr_0
    process(ptr_deref_2049_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2049_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2049_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2049_base_resize
    process(iNsTr_3_2046) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2046;
      ov := iv(6 downto 0);
      ptr_deref_2049_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2049_gather_scatter
    process(ptr_deref_2049_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2049_data_0;
      ov(15 downto 0) := iv;
      tmp12_2050 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2049_root_address_inst
    process(ptr_deref_2049_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2049_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2049_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2061_addr_0
    process(ptr_deref_2061_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2061_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2061_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2061_base_resize
    process(iNsTr_4_2058) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2058;
      ov := iv(6 downto 0);
      ptr_deref_2061_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2061_gather_scatter
    process(ptr_deref_2061_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2061_data_0;
      ov(15 downto 0) := iv;
      tmp16_2062 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2061_root_address_inst
    process(ptr_deref_2061_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2061_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2061_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2071_addr_0
    process(ptr_deref_2071_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2071_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2071_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2071_base_resize
    process(iNsTr_5_2068) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2068;
      ov := iv(0 downto 0);
      ptr_deref_2071_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2071_gather_scatter
    process(ptr_deref_2071_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2071_data_0;
      ov(15 downto 0) := iv;
      tmp25_2072 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2071_root_address_inst
    process(ptr_deref_2071_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2071_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2071_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2083_addr_0
    process(ptr_deref_2083_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2083_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2083_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2083_base_resize
    process(iNsTr_6_2080) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2080;
      ov := iv(6 downto 0);
      ptr_deref_2083_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2083_gather_scatter
    process(ptr_deref_2083_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2083_data_0;
      ov(15 downto 0) := iv;
      tmp28_2084 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2083_root_address_inst
    process(ptr_deref_2083_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2083_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2083_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2096_addr_0
    process(ptr_deref_2096_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2096_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2096_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2096_base_resize
    process(iNsTr_7_2093) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2093;
      ov := iv(0 downto 0);
      ptr_deref_2096_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2096_gather_scatter
    process(ptr_deref_2096_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2096_data_0;
      ov(15 downto 0) := iv;
      tmp37_2097 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2096_root_address_inst
    process(ptr_deref_2096_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2096_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2096_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2108_addr_0
    process(ptr_deref_2108_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2108_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2108_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2108_base_resize
    process(iNsTr_8_2105) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2105;
      ov := iv(6 downto 0);
      ptr_deref_2108_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2108_gather_scatter
    process(ptr_deref_2108_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2108_data_0;
      ov(15 downto 0) := iv;
      tmp40_2109 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2108_root_address_inst
    process(ptr_deref_2108_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2108_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2108_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2120_addr_0
    process(ptr_deref_2120_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2120_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2120_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2120_base_resize
    process(iNsTr_9_2117) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2117;
      ov := iv(6 downto 0);
      ptr_deref_2120_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2120_gather_scatter
    process(ptr_deref_2120_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2120_data_0;
      ov(15 downto 0) := iv;
      tmp50_2121 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2120_root_address_inst
    process(ptr_deref_2120_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2120_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2120_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2132_addr_0
    process(ptr_deref_2132_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2132_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2132_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2132_base_resize
    process(iNsTr_10_2129) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2129;
      ov := iv(6 downto 0);
      ptr_deref_2132_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2132_gather_scatter
    process(ptr_deref_2132_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2132_data_0;
      ov(15 downto 0) := iv;
      tmp54_2133 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2132_root_address_inst
    process(ptr_deref_2132_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2132_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2132_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2281_addr_0
    process(ptr_deref_2281_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2281_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2281_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2281_base_resize
    process(arrayidx_2278) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2278;
      ov := iv(13 downto 0);
      ptr_deref_2281_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2281_gather_scatter
    process(ptr_deref_2281_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2281_data_0;
      ov(63 downto 0) := iv;
      tmp65_2282 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2281_root_address_inst
    process(ptr_deref_2281_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2281_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2281_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2301_addr_0
    process(ptr_deref_2301_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2301_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2301_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2301_base_resize
    process(arrayidx70_2299) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx70_2299;
      ov := iv(13 downto 0);
      ptr_deref_2301_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2301_gather_scatter
    process(tmp65_2282) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp65_2282;
      ov(63 downto 0) := iv;
      ptr_deref_2301_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2301_root_address_inst
    process(ptr_deref_2301_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2301_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2301_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2319_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2318;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2319_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2319_branch_req_0,
          ack0 => if_stmt_2319_branch_ack_0,
          ack1 => if_stmt_2319_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2370_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp97_2369;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2370_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2370_branch_req_0,
          ack0 => if_stmt_2370_branch_ack_0,
          ack1 => if_stmt_2370_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2152_inst
    process(tmp40_2109) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp40_2109, type_cast_2151_wire_constant, tmp_var);
      tmp3_2153 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2163_inst
    process(tmp28_2084) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp28_2084, type_cast_2162_wire_constant, tmp_var);
      tmp7_2164 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2194_inst
    process(input_dim1x_x1x_xph_2172, tmp127_2190) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2172, tmp127_2190, tmp_var);
      tmp128_2195 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2209_inst
    process(tmp4_2158, tmp5_2205) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp4_2158, tmp5_2205, tmp_var);
      tmp6_2210 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2219_inst
    process(tmp8_2169, tmp9_2215) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp8_2169, tmp9_2215, tmp_var);
      tmp10_2220 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2229_inst
    process(tmp6_2210, tmp11_2225) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp6_2210, tmp11_2225, tmp_var);
      tmp13_2230 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2255_inst
    process(tmp129_2200, input_dim2x_x1_2251) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp129_2200, input_dim2x_x1_2251, tmp_var);
      add21_2256 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2260_inst
    process(tmp14_2235, input_dim2x_x1_2251) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_2235, input_dim2x_x1_2251, tmp_var);
      add61_2261 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2330_inst
    process(indvar_2238) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2238, type_cast_2329_wire_constant, tmp_var);
      indvarx_xnext_2331 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2338_inst
    process(input_dim1x_x1x_xph_2172) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2172, type_cast_2337_wire_constant, tmp_var);
      inc_2339 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2356_inst
    process(inc92_2352, input_dim0x_x2x_xph_2179) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc92_2352, input_dim0x_x2x_xph_2179, tmp_var);
      inc92x_xinput_dim0x_x2_2357 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2312_inst
    process(conv73_2307) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv73_2307, type_cast_2311_wire_constant, tmp_var);
      add74_2313 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2368_inst
    process(inc92x_xinput_dim0x_x2_2357, tmp_2032) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc92x_xinput_dim0x_x2_2357, tmp_2032, tmp_var);
      cmp97_2369 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2347_inst
    process(conv84_2343, div87_2147) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv84_2343, div87_2147, tmp_var);
      cmp88_2348 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2037_inst
    process(tmp_2032) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2032, type_cast_2036_wire_constant, tmp_var);
      div_2038 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2146_inst
    process(conv86_2141) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv86_2141, type_cast_2145_wire_constant, tmp_var);
      div87_2147 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2270_inst
    process(conv64_2265) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv64_2265, type_cast_2269_wire_constant, tmp_var);
      shr111_2271 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2291_inst
    process(conv67_2286) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv67_2286, type_cast_2290_wire_constant, tmp_var);
      shr68113_2292 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2189_inst
    process(tmp16_2062, input_dim0x_x2x_xph_2179) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_2062, input_dim0x_x2x_xph_2179, tmp_var);
      tmp127_2190 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2199_inst
    process(tmp12_2050, tmp128_2195) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_2050, tmp128_2195, tmp_var);
      tmp129_2200 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2204_inst
    process(tmp37_2097, input_dim1x_x1x_xph_2172) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp37_2097, input_dim1x_x1x_xph_2172, tmp_var);
      tmp5_2205 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2214_inst
    process(tmp25_2072, input_dim0x_x2x_xph_2179) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp25_2072, input_dim0x_x2x_xph_2179, tmp_var);
      tmp9_2215 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2224_inst
    process(tmp54_2133, tmp10_2220) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_2133, tmp10_2220, tmp_var);
      tmp11_2225 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2234_inst
    process(tmp50_2121, tmp13_2230) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp50_2121, tmp13_2230, tmp_var);
      tmp14_2235 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2250_inst
    process(indvar_2238) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2238, type_cast_2249_wire_constant, tmp_var);
      input_dim2x_x1_2251 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2157_inst
    process(tmp3_2153, tmp31_2087) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp3_2153, tmp31_2087, tmp_var);
      tmp4_2158 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2168_inst
    process(tmp7_2164, tmp31_2087) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp7_2164, tmp31_2087, tmp_var);
      tmp8_2169 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2317_inst
    process(add74_2313, conv76_2137) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add74_2313, conv76_2137, tmp_var);
      cmp_2318 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_2276_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr111_2275_scaled;
      array_obj_ref_2276_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2276_index_offset_req_0;
      array_obj_ref_2276_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2276_index_offset_req_1;
      array_obj_ref_2276_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_2297_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr68113_2296_scaled;
      array_obj_ref_2297_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2297_index_offset_req_0;
      array_obj_ref_2297_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2297_index_offset_req_1;
      array_obj_ref_2297_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : LOAD_padding_2086_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2086_load_0_req_0;
      LOAD_padding_2086_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2086_load_0_req_1;
      LOAD_padding_2086_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2086_word_address_0;
      LOAD_padding_2086_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2031_load_0 ptr_deref_2049_load_0 ptr_deref_2061_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2031_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2049_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2061_load_0_req_0;
      ptr_deref_2031_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2049_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2061_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2031_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2049_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2061_load_0_req_1;
      ptr_deref_2031_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2049_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2061_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2031_word_address_0 & ptr_deref_2049_word_address_0 & ptr_deref_2061_word_address_0;
      ptr_deref_2031_data_0 <= data_out(47 downto 32);
      ptr_deref_2049_data_0 <= data_out(31 downto 16);
      ptr_deref_2061_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2096_load_0 ptr_deref_2071_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2096_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2071_load_0_req_0;
      ptr_deref_2096_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2071_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2096_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2071_load_0_req_1;
      ptr_deref_2096_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2071_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2096_word_address_0 & ptr_deref_2071_word_address_0;
      ptr_deref_2096_data_0 <= data_out(31 downto 16);
      ptr_deref_2071_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2083_load_0 ptr_deref_2108_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2083_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2108_load_0_req_0;
      ptr_deref_2083_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2108_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2083_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2108_load_0_req_1;
      ptr_deref_2083_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2108_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2083_word_address_0 & ptr_deref_2108_word_address_0;
      ptr_deref_2083_data_0 <= data_out(31 downto 16);
      ptr_deref_2108_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2120_load_0 ptr_deref_2132_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2120_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2132_load_0_req_0;
      ptr_deref_2120_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2132_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2120_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2132_load_0_req_1;
      ptr_deref_2120_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2132_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2120_word_address_0 & ptr_deref_2132_word_address_0;
      ptr_deref_2120_data_0 <= data_out(31 downto 16);
      ptr_deref_2132_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2281_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2281_load_0_req_0;
      ptr_deref_2281_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2281_load_0_req_1;
      ptr_deref_2281_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2281_word_address_0;
      ptr_deref_2281_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2301_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2301_store_0_req_0;
      ptr_deref_2301_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2301_store_0_req_1;
      ptr_deref_2301_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2301_word_address_0;
      data_in <= ptr_deref_2301_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2018_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_start_2018_inst_req_0;
      RPIPE_Block2_start_2018_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_start_2018_inst_req_1;
      RPIPE_Block2_start_2018_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2019 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2378_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2378_inst_req_0;
      WPIPE_Block2_done_2378_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2378_inst_req_1;
      WPIPE_Block2_done_2378_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2019;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6990_start: Boolean;
  signal convTransposeD_CP_6990_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2437_load_0_ack_0 : boolean;
  signal ptr_deref_2437_load_0_req_1 : boolean;
  signal ptr_deref_2437_load_0_req_0 : boolean;
  signal ptr_deref_2437_load_0_ack_1 : boolean;
  signal ptr_deref_2419_load_0_req_0 : boolean;
  signal ptr_deref_2419_load_0_ack_0 : boolean;
  signal ptr_deref_2419_load_0_req_1 : boolean;
  signal ptr_deref_2419_load_0_ack_1 : boolean;
  signal RPIPE_Block3_start_2388_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2388_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2388_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2388_inst_ack_1 : boolean;
  signal ptr_deref_2401_load_0_req_0 : boolean;
  signal ptr_deref_2401_load_0_ack_0 : boolean;
  signal ptr_deref_2401_load_0_req_1 : boolean;
  signal ptr_deref_2401_load_0_ack_1 : boolean;
  signal ptr_deref_2447_load_0_req_0 : boolean;
  signal ptr_deref_2447_load_0_ack_0 : boolean;
  signal ptr_deref_2447_load_0_req_1 : boolean;
  signal ptr_deref_2447_load_0_ack_1 : boolean;
  signal ptr_deref_2459_load_0_req_0 : boolean;
  signal ptr_deref_2459_load_0_ack_0 : boolean;
  signal ptr_deref_2459_load_0_req_1 : boolean;
  signal ptr_deref_2459_load_0_ack_1 : boolean;
  signal LOAD_padding_2462_load_0_req_0 : boolean;
  signal LOAD_padding_2462_load_0_ack_0 : boolean;
  signal LOAD_padding_2462_load_0_req_1 : boolean;
  signal LOAD_padding_2462_load_0_ack_1 : boolean;
  signal ptr_deref_2472_load_0_req_0 : boolean;
  signal ptr_deref_2472_load_0_ack_0 : boolean;
  signal ptr_deref_2472_load_0_req_1 : boolean;
  signal ptr_deref_2472_load_0_ack_1 : boolean;
  signal ptr_deref_2484_load_0_req_0 : boolean;
  signal ptr_deref_2484_load_0_ack_0 : boolean;
  signal ptr_deref_2484_load_0_req_1 : boolean;
  signal ptr_deref_2484_load_0_ack_1 : boolean;
  signal ptr_deref_2496_load_0_req_0 : boolean;
  signal ptr_deref_2496_load_0_ack_0 : boolean;
  signal ptr_deref_2496_load_0_req_1 : boolean;
  signal ptr_deref_2496_load_0_ack_1 : boolean;
  signal ptr_deref_2508_load_0_req_0 : boolean;
  signal ptr_deref_2508_load_0_ack_0 : boolean;
  signal ptr_deref_2508_load_0_req_1 : boolean;
  signal ptr_deref_2508_load_0_ack_1 : boolean;
  signal type_cast_2512_inst_req_0 : boolean;
  signal type_cast_2512_inst_ack_0 : boolean;
  signal type_cast_2512_inst_req_1 : boolean;
  signal type_cast_2512_inst_ack_1 : boolean;
  signal type_cast_2629_inst_req_0 : boolean;
  signal type_cast_2629_inst_ack_0 : boolean;
  signal type_cast_2629_inst_req_1 : boolean;
  signal type_cast_2629_inst_ack_1 : boolean;
  signal array_obj_ref_2641_index_offset_req_0 : boolean;
  signal array_obj_ref_2641_index_offset_ack_0 : boolean;
  signal array_obj_ref_2641_index_offset_req_1 : boolean;
  signal array_obj_ref_2641_index_offset_ack_1 : boolean;
  signal addr_of_2642_final_reg_req_0 : boolean;
  signal addr_of_2642_final_reg_ack_0 : boolean;
  signal addr_of_2642_final_reg_req_1 : boolean;
  signal addr_of_2642_final_reg_ack_1 : boolean;
  signal ptr_deref_2646_load_0_req_0 : boolean;
  signal ptr_deref_2646_load_0_ack_0 : boolean;
  signal ptr_deref_2646_load_0_req_1 : boolean;
  signal ptr_deref_2646_load_0_ack_1 : boolean;
  signal type_cast_2650_inst_req_0 : boolean;
  signal type_cast_2650_inst_ack_0 : boolean;
  signal type_cast_2650_inst_req_1 : boolean;
  signal type_cast_2650_inst_ack_1 : boolean;
  signal array_obj_ref_2662_index_offset_req_0 : boolean;
  signal array_obj_ref_2662_index_offset_ack_0 : boolean;
  signal array_obj_ref_2662_index_offset_req_1 : boolean;
  signal array_obj_ref_2662_index_offset_ack_1 : boolean;
  signal addr_of_2663_final_reg_req_0 : boolean;
  signal addr_of_2663_final_reg_ack_0 : boolean;
  signal addr_of_2663_final_reg_req_1 : boolean;
  signal addr_of_2663_final_reg_ack_1 : boolean;
  signal ptr_deref_2666_store_0_req_0 : boolean;
  signal ptr_deref_2666_store_0_ack_0 : boolean;
  signal ptr_deref_2666_store_0_req_1 : boolean;
  signal ptr_deref_2666_store_0_ack_1 : boolean;
  signal type_cast_2671_inst_req_0 : boolean;
  signal type_cast_2671_inst_ack_0 : boolean;
  signal type_cast_2671_inst_req_1 : boolean;
  signal type_cast_2671_inst_ack_1 : boolean;
  signal if_stmt_2684_branch_req_0 : boolean;
  signal if_stmt_2684_branch_ack_1 : boolean;
  signal if_stmt_2684_branch_ack_0 : boolean;
  signal if_stmt_2739_branch_req_0 : boolean;
  signal if_stmt_2739_branch_ack_1 : boolean;
  signal if_stmt_2739_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2747_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2747_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2747_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2747_inst_ack_1 : boolean;
  signal type_cast_2543_inst_req_0 : boolean;
  signal type_cast_2543_inst_ack_0 : boolean;
  signal type_cast_2543_inst_req_1 : boolean;
  signal type_cast_2543_inst_ack_1 : boolean;
  signal phi_stmt_2538_req_1 : boolean;
  signal type_cast_2547_inst_req_0 : boolean;
  signal type_cast_2547_inst_ack_0 : boolean;
  signal type_cast_2547_inst_req_1 : boolean;
  signal type_cast_2547_inst_ack_1 : boolean;
  signal phi_stmt_2544_req_0 : boolean;
  signal type_cast_2541_inst_req_0 : boolean;
  signal type_cast_2541_inst_ack_0 : boolean;
  signal type_cast_2541_inst_req_1 : boolean;
  signal type_cast_2541_inst_ack_1 : boolean;
  signal phi_stmt_2538_req_0 : boolean;
  signal type_cast_2549_inst_req_0 : boolean;
  signal type_cast_2549_inst_ack_0 : boolean;
  signal type_cast_2549_inst_req_1 : boolean;
  signal type_cast_2549_inst_ack_1 : boolean;
  signal phi_stmt_2544_req_1 : boolean;
  signal phi_stmt_2538_ack_0 : boolean;
  signal phi_stmt_2544_ack_0 : boolean;
  signal type_cast_2609_inst_req_0 : boolean;
  signal type_cast_2609_inst_ack_0 : boolean;
  signal type_cast_2609_inst_req_1 : boolean;
  signal type_cast_2609_inst_ack_1 : boolean;
  signal phi_stmt_2603_req_1 : boolean;
  signal phi_stmt_2603_req_0 : boolean;
  signal phi_stmt_2603_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6990_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6990_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6990_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6990_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6990: Block -- control-path 
    signal convTransposeD_CP_6990_elements: BooleanArray(75 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6990_elements(0) <= convTransposeD_CP_6990_start;
    convTransposeD_CP_6990_symbol <= convTransposeD_CP_6990_elements(51);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2386/$entry
      -- CP-element group 0: 	 branch_block_stmt_2386/branch_block_stmt_2386__entry__
      -- CP-element group 0: 	 branch_block_stmt_2386/assign_stmt_2389__entry__
      -- CP-element group 0: 	 branch_block_stmt_2386/assign_stmt_2389/$entry
      -- CP-element group 0: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_Sample/rr
      -- 
    rr_7038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(0), ack => RPIPE_Block3_start_2388_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_Update/cr
      -- 
    ra_7039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2388_inst_ack_0, ack => convTransposeD_CP_6990_elements(1)); -- 
    cr_7043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(1), ack => RPIPE_Block3_start_2388_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (256) 
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2389__exit__
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535__entry__
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2389/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2389/RPIPE_Block3_start_2388_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_Update/cr
      -- 
    ca_7044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2388_inst_ack_1, ack => convTransposeD_CP_6990_elements(2)); -- 
    cr_7191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2437_load_0_req_1); -- 
    rr_7180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2437_load_0_req_0); -- 
    rr_7130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2419_load_0_req_0); -- 
    cr_7141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2419_load_0_req_1); -- 
    rr_7080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2401_load_0_req_0); -- 
    cr_7091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2401_load_0_req_1); -- 
    rr_7230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2447_load_0_req_0); -- 
    cr_7241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2447_load_0_req_1); -- 
    rr_7280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2459_load_0_req_0); -- 
    cr_7291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2459_load_0_req_1); -- 
    rr_7313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => LOAD_padding_2462_load_0_req_0); -- 
    cr_7324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => LOAD_padding_2462_load_0_req_1); -- 
    rr_7363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2472_load_0_req_0); -- 
    cr_7374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2472_load_0_req_1); -- 
    rr_7413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2484_load_0_req_0); -- 
    cr_7424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2484_load_0_req_1); -- 
    rr_7463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2496_load_0_req_0); -- 
    cr_7474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2496_load_0_req_1); -- 
    rr_7513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2508_load_0_req_0); -- 
    cr_7524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => ptr_deref_2508_load_0_req_1); -- 
    cr_7543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(2), ack => type_cast_2512_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Sample/word_access_start/word_0/ra
      -- 
    ra_7081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2401_load_0_ack_0, ack => convTransposeD_CP_6990_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	25 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/ptr_deref_2401_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/ptr_deref_2401_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/ptr_deref_2401_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2401_Update/ptr_deref_2401_Merge/merge_ack
      -- 
    ca_7092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2401_load_0_ack_1, ack => convTransposeD_CP_6990_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_sample_completed_
      -- 
    ra_7131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2419_load_0_ack_0, ack => convTransposeD_CP_6990_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	25 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/ptr_deref_2419_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/ptr_deref_2419_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/ptr_deref_2419_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2419_Update/ptr_deref_2419_Merge/$entry
      -- 
    ca_7142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2419_load_0_ack_1, ack => convTransposeD_CP_6990_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Sample/$exit
      -- 
    ra_7181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2437_load_0_ack_0, ack => convTransposeD_CP_6990_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/ptr_deref_2437_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/ptr_deref_2437_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/ptr_deref_2437_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/ptr_deref_2437_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2437_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_Sample/rr
      -- 
    ca_7192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2437_load_0_ack_1, ack => convTransposeD_CP_6990_elements(8)); -- 
    rr_7538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(8), ack => type_cast_2512_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Sample/word_access_start/word_0/ra
      -- 
    ra_7231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2447_load_0_ack_0, ack => convTransposeD_CP_6990_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	25 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/ptr_deref_2447_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/ptr_deref_2447_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/ptr_deref_2447_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2447_Update/ptr_deref_2447_Merge/merge_ack
      -- 
    ca_7242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2447_load_0_ack_1, ack => convTransposeD_CP_6990_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Sample/word_access_start/word_0/ra
      -- 
    ra_7281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2459_load_0_ack_0, ack => convTransposeD_CP_6990_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	25 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/ptr_deref_2459_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/ptr_deref_2459_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/ptr_deref_2459_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2459_Update/ptr_deref_2459_Merge/merge_ack
      -- 
    ca_7292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2459_load_0_ack_1, ack => convTransposeD_CP_6990_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Sample/word_access_start/word_0/ra
      -- 
    ra_7314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2462_load_0_ack_0, ack => convTransposeD_CP_6990_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	25 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/LOAD_padding_2462_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/LOAD_padding_2462_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/LOAD_padding_2462_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/LOAD_padding_2462_Update/LOAD_padding_2462_Merge/merge_ack
      -- 
    ca_7325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2462_load_0_ack_1, ack => convTransposeD_CP_6990_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Sample/word_access_start/word_0/ra
      -- 
    ra_7364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2472_load_0_ack_0, ack => convTransposeD_CP_6990_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	25 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/ptr_deref_2472_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/ptr_deref_2472_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/ptr_deref_2472_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2472_Update/ptr_deref_2472_Merge/merge_ack
      -- 
    ca_7375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2472_load_0_ack_1, ack => convTransposeD_CP_6990_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Sample/word_access_start/word_0/ra
      -- 
    ra_7414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2484_load_0_ack_0, ack => convTransposeD_CP_6990_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/ptr_deref_2484_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/ptr_deref_2484_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/ptr_deref_2484_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2484_Update/ptr_deref_2484_Merge/merge_ack
      -- 
    ca_7425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2484_load_0_ack_1, ack => convTransposeD_CP_6990_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Sample/word_access_start/word_0/ra
      -- 
    ra_7464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2496_load_0_ack_0, ack => convTransposeD_CP_6990_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	25 
    -- CP-element group 20:  members (9) 
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/ptr_deref_2496_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/ptr_deref_2496_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/ptr_deref_2496_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2496_Update/ptr_deref_2496_Merge/merge_ack
      -- 
    ca_7475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2496_load_0_ack_1, ack => convTransposeD_CP_6990_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Sample/word_access_start/word_0/ra
      -- 
    ra_7514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2508_load_0_ack_0, ack => convTransposeD_CP_6990_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/ptr_deref_2508_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/ptr_deref_2508_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/ptr_deref_2508_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/ptr_deref_2508_Update/ptr_deref_2508_Merge/merge_ack
      -- 
    ca_7525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2508_load_0_ack_1, ack => convTransposeD_CP_6990_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_Sample/ra
      -- 
    ra_7539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_0, ack => convTransposeD_CP_6990_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/type_cast_2512_Update/ca
      -- 
    ca_7544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2512_inst_ack_1, ack => convTransposeD_CP_6990_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  place  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: 	18 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	22 
    -- CP-element group 25: 	16 
    -- CP-element group 25: 	14 
    -- CP-element group 25: 	4 
    -- CP-element group 25: 	6 
    -- CP-element group 25: 	10 
    -- CP-element group 25: 	12 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	52 
    -- CP-element group 25: 	53 
    -- CP-element group 25: 	55 
    -- CP-element group 25: 	56 
    -- CP-element group 25:  members (20) 
      -- CP-element group 25: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535__exit__
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter
      -- CP-element group 25: 	 branch_block_stmt_2386/assign_stmt_2398_to_assign_stmt_2535/$exit
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/Update/cr
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/Update/cr
      -- 
    rr_7864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(25), ack => type_cast_2543_inst_req_0); -- 
    cr_7869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(25), ack => type_cast_2543_inst_req_1); -- 
    rr_7887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(25), ack => type_cast_2547_inst_req_0); -- 
    cr_7892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(25), ack => type_cast_2547_inst_req_1); -- 
    convTransposeD_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(24) & convTransposeD_CP_6990_elements(18) & convTransposeD_CP_6990_elements(20) & convTransposeD_CP_6990_elements(22) & convTransposeD_CP_6990_elements(16) & convTransposeD_CP_6990_elements(14) & convTransposeD_CP_6990_elements(4) & convTransposeD_CP_6990_elements(6) & convTransposeD_CP_6990_elements(10) & convTransposeD_CP_6990_elements(12);
      gj_convTransposeD_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	75 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_Sample/ra
      -- 
    ra_7559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2629_inst_ack_0, ack => convTransposeD_CP_6990_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	75 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (16) 
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_resize_1/index_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_Sample/req
      -- 
    ca_7564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2629_inst_ack_1, ack => convTransposeD_CP_6990_elements(27)); -- 
    req_7589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(27), ack => array_obj_ref_2641_index_offset_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	45 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_sample_complete
      -- CP-element group 28: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_Sample/ack
      -- 
    ack_7590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2641_index_offset_ack_0, ack => convTransposeD_CP_6990_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	75 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (11) 
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_root_address_calculated
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_offset_calculated
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_Update/ack
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_base_plus_offset/$entry
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_base_plus_offset/$exit
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_base_plus_offset/sum_rename_req
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_base_plus_offset/sum_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_request/$entry
      -- CP-element group 29: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_request/req
      -- 
    ack_7595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2641_index_offset_ack_1, ack => convTransposeD_CP_6990_elements(29)); -- 
    req_7604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(29), ack => addr_of_2642_final_reg_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_request/$exit
      -- CP-element group 30: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_request/ack
      -- 
    ack_7605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2642_final_reg_ack_0, ack => convTransposeD_CP_6990_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	75 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (24) 
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_complete/$exit
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_complete/ack
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_word_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_root_address_calculated
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_address_resized
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_addr_resize/$entry
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_addr_resize/$exit
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_addr_resize/base_resize_req
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_addr_resize/base_resize_ack
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_plus_offset/$entry
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_plus_offset/$exit
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_plus_offset/sum_rename_req
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_base_plus_offset/sum_rename_ack
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_word_addrgen/$entry
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_word_addrgen/$exit
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_word_addrgen/root_register_req
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_word_addrgen/root_register_ack
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Sample/word_access_start/word_0/rr
      -- 
    ack_7610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2642_final_reg_ack_1, ack => convTransposeD_CP_6990_elements(31)); -- 
    rr_7643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(31), ack => ptr_deref_2646_load_0_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Sample/word_access_start/$exit
      -- CP-element group 32: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Sample/word_access_start/word_0/ra
      -- 
    ra_7644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2646_load_0_ack_0, ack => convTransposeD_CP_6990_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	75 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	40 
    -- CP-element group 33:  members (9) 
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/word_access_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/word_access_complete/word_0/ca
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/ptr_deref_2646_Merge/$entry
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/ptr_deref_2646_Merge/$exit
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/ptr_deref_2646_Merge/merge_req
      -- CP-element group 33: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/ptr_deref_2646_Merge/merge_ack
      -- 
    ca_7655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2646_load_0_ack_1, ack => convTransposeD_CP_6990_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	75 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_Sample/ra
      -- 
    ra_7669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2650_inst_ack_0, ack => convTransposeD_CP_6990_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	75 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_Sample/req
      -- 
    ca_7674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2650_inst_ack_1, ack => convTransposeD_CP_6990_elements(35)); -- 
    req_7699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(35), ack => array_obj_ref_2662_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	45 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_Sample/ack
      -- 
    ack_7700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2662_index_offset_ack_0, ack => convTransposeD_CP_6990_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	75 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_request/req
      -- 
    ack_7705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2662_index_offset_ack_1, ack => convTransposeD_CP_6990_elements(37)); -- 
    req_7714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(37), ack => addr_of_2663_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_request/ack
      -- 
    ack_7715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2663_final_reg_ack_0, ack => convTransposeD_CP_6990_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	75 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (19) 
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_word_addrgen/root_register_ack
      -- 
    ack_7720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2663_final_reg_ack_1, ack => convTransposeD_CP_6990_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	33 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/ptr_deref_2666_Split/$entry
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/ptr_deref_2666_Split/$exit
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/ptr_deref_2666_Split/split_req
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/ptr_deref_2666_Split/split_ack
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/word_access_start/$entry
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/word_access_start/word_0/$entry
      -- CP-element group 40: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/word_access_start/word_0/rr
      -- 
    rr_7758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(40), ack => ptr_deref_2666_store_0_req_0); -- 
    convTransposeD_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(33) & convTransposeD_CP_6990_elements(39);
      gj_convTransposeD_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/word_access_start/$exit
      -- CP-element group 41: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/word_access_start/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Sample/word_access_start/word_0/ra
      -- 
    ra_7759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2666_store_0_ack_0, ack => convTransposeD_CP_6990_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	75 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Update/word_access_complete/$exit
      -- CP-element group 42: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Update/word_access_complete/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Update/word_access_complete/word_0/ca
      -- 
    ca_7770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2666_store_0_ack_1, ack => convTransposeD_CP_6990_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	75 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_Sample/ra
      -- 
    ra_7779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2671_inst_ack_0, ack => convTransposeD_CP_6990_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	75 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_Update/ca
      -- 
    ca_7784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2671_inst_ack_1, ack => convTransposeD_CP_6990_elements(44)); -- 
    -- CP-element group 45:  branch  join  transition  place  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	28 
    -- CP-element group 45: 	36 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (10) 
      -- CP-element group 45: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683__exit__
      -- CP-element group 45: 	 branch_block_stmt_2386/if_stmt_2684__entry__
      -- CP-element group 45: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/$exit
      -- CP-element group 45: 	 branch_block_stmt_2386/if_stmt_2684_dead_link/$entry
      -- CP-element group 45: 	 branch_block_stmt_2386/if_stmt_2684_eval_test/$entry
      -- CP-element group 45: 	 branch_block_stmt_2386/if_stmt_2684_eval_test/$exit
      -- CP-element group 45: 	 branch_block_stmt_2386/if_stmt_2684_eval_test/branch_req
      -- CP-element group 45: 	 branch_block_stmt_2386/R_cmp_2685_place
      -- CP-element group 45: 	 branch_block_stmt_2386/if_stmt_2684_if_link/$entry
      -- CP-element group 45: 	 branch_block_stmt_2386/if_stmt_2684_else_link/$entry
      -- 
    branch_req_7792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(45), ack => if_stmt_2684_branch_req_0); -- 
    convTransposeD_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(42) & convTransposeD_CP_6990_elements(44) & convTransposeD_CP_6990_elements(28) & convTransposeD_CP_6990_elements(36);
      gj_convTransposeD_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	70 
    -- CP-element group 46: 	71 
    -- CP-element group 46:  members (24) 
      -- CP-element group 46: 	 branch_block_stmt_2386/merge_stmt_2690_PhiAck/$exit
      -- CP-element group 46: 	 branch_block_stmt_2386/merge_stmt_2690_PhiAck/dummy
      -- CP-element group 46: 	 branch_block_stmt_2386/merge_stmt_2690_PhiAck/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/merge_stmt_2690__exit__
      -- CP-element group 46: 	 branch_block_stmt_2386/assign_stmt_2696__entry__
      -- CP-element group 46: 	 branch_block_stmt_2386/assign_stmt_2696__exit__
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody
      -- CP-element group 46: 	 branch_block_stmt_2386/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 46: 	 branch_block_stmt_2386/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/merge_stmt_2690_PhiReqMerge
      -- CP-element group 46: 	 branch_block_stmt_2386/if_stmt_2684_if_link/$exit
      -- CP-element group 46: 	 branch_block_stmt_2386/if_stmt_2684_if_link/if_choice_transition
      -- CP-element group 46: 	 branch_block_stmt_2386/whilex_xbody_ifx_xthen
      -- CP-element group 46: 	 branch_block_stmt_2386/assign_stmt_2696/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/assign_stmt_2696/$exit
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2684_branch_ack_1, ack => convTransposeD_CP_6990_elements(46)); -- 
    rr_7968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(46), ack => type_cast_2609_inst_req_0); -- 
    cr_7973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(46), ack => type_cast_2609_inst_req_1); -- 
    -- CP-element group 47:  branch  transition  place  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (22) 
      -- CP-element group 47: 	 branch_block_stmt_2386/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 47: 	 branch_block_stmt_2386/merge_stmt_2698_PhiReqMerge
      -- CP-element group 47: 	 branch_block_stmt_2386/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 47: 	 branch_block_stmt_2386/merge_stmt_2698__exit__
      -- CP-element group 47: 	 branch_block_stmt_2386/assign_stmt_2704_to_assign_stmt_2738__entry__
      -- CP-element group 47: 	 branch_block_stmt_2386/assign_stmt_2704_to_assign_stmt_2738__exit__
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2739__entry__
      -- CP-element group 47: 	 branch_block_stmt_2386/merge_stmt_2698_PhiAck/dummy
      -- CP-element group 47: 	 branch_block_stmt_2386/merge_stmt_2698_PhiAck/$exit
      -- CP-element group 47: 	 branch_block_stmt_2386/merge_stmt_2698_PhiAck/$entry
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2684_else_link/$exit
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2684_else_link/else_choice_transition
      -- CP-element group 47: 	 branch_block_stmt_2386/whilex_xbody_ifx_xelse
      -- CP-element group 47: 	 branch_block_stmt_2386/assign_stmt_2704_to_assign_stmt_2738/$entry
      -- CP-element group 47: 	 branch_block_stmt_2386/assign_stmt_2704_to_assign_stmt_2738/$exit
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2739_dead_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2739_eval_test/$entry
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2739_eval_test/$exit
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2739_eval_test/branch_req
      -- CP-element group 47: 	 branch_block_stmt_2386/R_cmp104_2740_place
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2739_if_link/$entry
      -- CP-element group 47: 	 branch_block_stmt_2386/if_stmt_2739_else_link/$entry
      -- 
    else_choice_transition_7801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2684_branch_ack_0, ack => convTransposeD_CP_6990_elements(47)); -- 
    branch_req_7817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(47), ack => if_stmt_2739_branch_req_0); -- 
    -- CP-element group 48:  merge  transition  place  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (15) 
      -- CP-element group 48: 	 branch_block_stmt_2386/merge_stmt_2745_PhiAck/$entry
      -- CP-element group 48: 	 branch_block_stmt_2386/merge_stmt_2745_PhiReqMerge
      -- CP-element group 48: 	 branch_block_stmt_2386/merge_stmt_2745_PhiAck/$exit
      -- CP-element group 48: 	 branch_block_stmt_2386/merge_stmt_2745_PhiAck/dummy
      -- CP-element group 48: 	 branch_block_stmt_2386/merge_stmt_2745__exit__
      -- CP-element group 48: 	 branch_block_stmt_2386/assign_stmt_2749__entry__
      -- CP-element group 48: 	 branch_block_stmt_2386/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 48: 	 branch_block_stmt_2386/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 48: 	 branch_block_stmt_2386/if_stmt_2739_if_link/$exit
      -- CP-element group 48: 	 branch_block_stmt_2386/if_stmt_2739_if_link/if_choice_transition
      -- CP-element group 48: 	 branch_block_stmt_2386/ifx_xelse_whilex_xend
      -- CP-element group 48: 	 branch_block_stmt_2386/assign_stmt_2749/$entry
      -- CP-element group 48: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_Sample/req
      -- 
    if_choice_transition_7822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2739_branch_ack_1, ack => convTransposeD_CP_6990_elements(48)); -- 
    req_7839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(48), ack => WPIPE_Block3_done_2747_inst_req_0); -- 
    -- CP-element group 49:  fork  transition  place  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	62 
    -- CP-element group 49: 	63 
    -- CP-element group 49: 	60 
    -- CP-element group 49: 	59 
    -- CP-element group 49:  members (20) 
      -- CP-element group 49: 	 branch_block_stmt_2386/if_stmt_2739_else_link/$exit
      -- CP-element group 49: 	 branch_block_stmt_2386/if_stmt_2739_else_link/else_choice_transition
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/Update/cr
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/Sample/rr
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2739_branch_ack_0, ack => convTransposeD_CP_6990_elements(49)); -- 
    rr_7913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(49), ack => type_cast_2541_inst_req_0); -- 
    cr_7918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(49), ack => type_cast_2541_inst_req_1); -- 
    rr_7936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(49), ack => type_cast_2549_inst_req_0); -- 
    cr_7941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(49), ack => type_cast_2549_inst_req_1); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_update_start_
      -- CP-element group 50: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_Update/req
      -- 
    ack_7840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2747_inst_ack_0, ack => convTransposeD_CP_6990_elements(50)); -- 
    req_7844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(50), ack => WPIPE_Block3_done_2747_inst_req_1); -- 
    -- CP-element group 51:  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2386/merge_stmt_2751_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_2386/return___PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_2386/return___PhiReq/$exit
      -- CP-element group 51: 	 $exit
      -- CP-element group 51: 	 branch_block_stmt_2386/$exit
      -- CP-element group 51: 	 branch_block_stmt_2386/branch_block_stmt_2386__exit__
      -- CP-element group 51: 	 branch_block_stmt_2386/assign_stmt_2749__exit__
      -- CP-element group 51: 	 branch_block_stmt_2386/return__
      -- CP-element group 51: 	 branch_block_stmt_2386/merge_stmt_2751__exit__
      -- CP-element group 51: 	 branch_block_stmt_2386/merge_stmt_2751_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_2386/merge_stmt_2751_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_2386/merge_stmt_2751_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_2386/assign_stmt_2749/$exit
      -- CP-element group 51: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2386/assign_stmt_2749/WPIPE_Block3_done_2747_Update/ack
      -- 
    ack_7845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2747_inst_ack_1, ack => convTransposeD_CP_6990_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	25 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/Sample/ra
      -- 
    ra_7865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2543_inst_ack_0, ack => convTransposeD_CP_6990_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	25 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/Update/ca
      -- 
    ca_7870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2543_inst_ack_1, ack => convTransposeD_CP_6990_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	58 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/$exit
      -- CP-element group 54: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/$exit
      -- CP-element group 54: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/$exit
      -- CP-element group 54: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2543/SplitProtocol/$exit
      -- CP-element group 54: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_req
      -- 
    phi_stmt_2538_req_7871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2538_req_7871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(54), ack => phi_stmt_2538_req_1); -- 
    convTransposeD_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(52) & convTransposeD_CP_6990_elements(53);
      gj_convTransposeD_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	25 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/Sample/ra
      -- 
    ra_7888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2547_inst_ack_0, ack => convTransposeD_CP_6990_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	25 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/Update/ca
      -- 
    ca_7893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2547_inst_ack_1, ack => convTransposeD_CP_6990_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/$exit
      -- CP-element group 57: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/$exit
      -- CP-element group 57: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/$exit
      -- CP-element group 57: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2547/SplitProtocol/$exit
      -- CP-element group 57: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_req
      -- 
    phi_stmt_2544_req_7894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2544_req_7894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(57), ack => phi_stmt_2544_req_0); -- 
    convTransposeD_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(55) & convTransposeD_CP_6990_elements(56);
      gj_convTransposeD_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	54 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	66 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_2386/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(54) & convTransposeD_CP_6990_elements(57);
      gj_convTransposeD_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	49 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/Sample/ra
      -- 
    ra_7914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2541_inst_ack_0, ack => convTransposeD_CP_6990_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	49 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/Update/ca
      -- 
    ca_7919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2541_inst_ack_1, ack => convTransposeD_CP_6990_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	65 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/$exit
      -- CP-element group 61: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/$exit
      -- CP-element group 61: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/$exit
      -- CP-element group 61: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_sources/type_cast_2541/SplitProtocol/$exit
      -- CP-element group 61: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2538/phi_stmt_2538_req
      -- 
    phi_stmt_2538_req_7920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2538_req_7920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(61), ack => phi_stmt_2538_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(60) & convTransposeD_CP_6990_elements(59);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	49 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/Sample/ra
      -- 
    ra_7937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2549_inst_ack_0, ack => convTransposeD_CP_6990_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	49 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/Update/ca
      -- 
    ca_7942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2549_inst_ack_1, ack => convTransposeD_CP_6990_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/$exit
      -- CP-element group 64: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/$exit
      -- CP-element group 64: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/$exit
      -- CP-element group 64: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_sources/type_cast_2549/SplitProtocol/$exit
      -- CP-element group 64: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2544/phi_stmt_2544_req
      -- 
    phi_stmt_2544_req_7943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2544_req_7943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(64), ack => phi_stmt_2544_req_1); -- 
    convTransposeD_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(62) & convTransposeD_CP_6990_elements(63);
      gj_convTransposeD_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: 	61 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_2386/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(64) & convTransposeD_CP_6990_elements(61);
      gj_convTransposeD_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  merge  fork  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: 	58 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_2386/merge_stmt_2537_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_2386/merge_stmt_2537_PhiAck/$entry
      -- 
    convTransposeD_CP_6990_elements(66) <= OrReduce(convTransposeD_CP_6990_elements(65) & convTransposeD_CP_6990_elements(58));
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_2386/merge_stmt_2537_PhiAck/phi_stmt_2538_ack
      -- 
    phi_stmt_2538_ack_7948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2538_ack_0, ack => convTransposeD_CP_6990_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_2386/merge_stmt_2537_PhiAck/phi_stmt_2544_ack
      -- 
    phi_stmt_2544_ack_7949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2544_ack_0, ack => convTransposeD_CP_6990_elements(68)); -- 
    -- CP-element group 69:  join  transition  place  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	73 
    -- CP-element group 69:  members (10) 
      -- CP-element group 69: 	 branch_block_stmt_2386/merge_stmt_2537__exit__
      -- CP-element group 69: 	 branch_block_stmt_2386/assign_stmt_2555_to_assign_stmt_2600__entry__
      -- CP-element group 69: 	 branch_block_stmt_2386/assign_stmt_2555_to_assign_stmt_2600__exit__
      -- CP-element group 69: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 69: 	 branch_block_stmt_2386/assign_stmt_2555_to_assign_stmt_2600/$entry
      -- CP-element group 69: 	 branch_block_stmt_2386/assign_stmt_2555_to_assign_stmt_2600/$exit
      -- CP-element group 69: 	 branch_block_stmt_2386/merge_stmt_2537_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2603/$entry
      -- CP-element group 69: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/$entry
      -- 
    convTransposeD_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(67) & convTransposeD_CP_6990_elements(68);
      gj_convTransposeD_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	46 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/Sample/ra
      -- 
    ra_7969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_0, ack => convTransposeD_CP_6990_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	46 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/Update/ca
      -- 
    ca_7974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2609_inst_ack_1, ack => convTransposeD_CP_6990_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/$exit
      -- CP-element group 72: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/$exit
      -- CP-element group 72: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/$exit
      -- CP-element group 72: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2609/SplitProtocol/$exit
      -- CP-element group 72: 	 branch_block_stmt_2386/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_req
      -- 
    phi_stmt_2603_req_7975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2603_req_7975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(72), ack => phi_stmt_2603_req_1); -- 
    convTransposeD_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6990_elements(70) & convTransposeD_CP_6990_elements(71);
      gj_convTransposeD_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6990_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  output  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 73: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2603/$exit
      -- CP-element group 73: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_sources/type_cast_2607_konst_delay_trans
      -- CP-element group 73: 	 branch_block_stmt_2386/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2603/phi_stmt_2603_req
      -- 
    phi_stmt_2603_req_7986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2603_req_7986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(73), ack => phi_stmt_2603_req_0); -- 
    -- Element group convTransposeD_CP_6990_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => convTransposeD_CP_6990_elements(69), ack => convTransposeD_CP_6990_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  merge  transition  place  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2386/merge_stmt_2602_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2386/merge_stmt_2602_PhiAck/$entry
      -- 
    convTransposeD_CP_6990_elements(74) <= OrReduce(convTransposeD_CP_6990_elements(72) & convTransposeD_CP_6990_elements(73));
    -- CP-element group 75:  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	34 
    -- CP-element group 75: 	42 
    -- CP-element group 75: 	43 
    -- CP-element group 75: 	44 
    -- CP-element group 75: 	33 
    -- CP-element group 75: 	31 
    -- CP-element group 75: 	26 
    -- CP-element group 75: 	37 
    -- CP-element group 75: 	27 
    -- CP-element group 75: 	29 
    -- CP-element group 75: 	35 
    -- CP-element group 75: 	39 
    -- CP-element group 75:  members (45) 
      -- CP-element group 75: 	 branch_block_stmt_2386/merge_stmt_2602__exit__
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683__entry__
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2629_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_update_start
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2641_final_index_sum_regn_Update/req
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2642_complete/req
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/word_access_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2646_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2650_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_update_start
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/array_obj_ref_2662_final_index_sum_regn_Update/req
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/addr_of_2663_complete/req
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Update/word_access_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/ptr_deref_2666_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2386/assign_stmt_2616_to_assign_stmt_2683/type_cast_2671_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_2386/merge_stmt_2602_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2386/merge_stmt_2602_PhiAck/phi_stmt_2603_ack
      -- 
    phi_stmt_2603_ack_7991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2603_ack_0, ack => convTransposeD_CP_6990_elements(75)); -- 
    rr_7558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => type_cast_2629_inst_req_0); -- 
    cr_7563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => type_cast_2629_inst_req_1); -- 
    req_7594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => array_obj_ref_2641_index_offset_req_1); -- 
    req_7609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => addr_of_2642_final_reg_req_1); -- 
    cr_7654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => ptr_deref_2646_load_0_req_1); -- 
    rr_7668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => type_cast_2650_inst_req_0); -- 
    cr_7673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => type_cast_2650_inst_req_1); -- 
    req_7704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => array_obj_ref_2662_index_offset_req_1); -- 
    req_7719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => addr_of_2663_final_reg_req_1); -- 
    cr_7769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => ptr_deref_2666_store_0_req_1); -- 
    rr_7778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => type_cast_2671_inst_req_0); -- 
    cr_7783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6990_elements(75), ack => type_cast_2671_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_padding_2462_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2462_word_address_0 : std_logic_vector(0 downto 0);
    signal R_shr118_2640_resized : std_logic_vector(13 downto 0);
    signal R_shr118_2640_scaled : std_logic_vector(13 downto 0);
    signal R_shr72120_2661_resized : std_logic_vector(13 downto 0);
    signal R_shr72120_2661_scaled : std_logic_vector(13 downto 0);
    signal add25_2621 : std_logic_vector(15 downto 0);
    signal add65_2626 : std_logic_vector(15 downto 0);
    signal add78_2678 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2641_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2641_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2641_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2641_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2641_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2641_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2662_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2662_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2662_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2662_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2662_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2662_root_address : std_logic_vector(13 downto 0);
    signal arrayidx74_2664 : std_logic_vector(31 downto 0);
    signal arrayidx_2643 : std_logic_vector(31 downto 0);
    signal call_2389 : std_logic_vector(15 downto 0);
    signal cmp104_2738 : std_logic_vector(0 downto 0);
    signal cmp91_2709 : std_logic_vector(0 downto 0);
    signal cmp_2683 : std_logic_vector(0 downto 0);
    signal conv68_2630 : std_logic_vector(63 downto 0);
    signal conv71_2651 : std_logic_vector(63 downto 0);
    signal conv77_2672 : std_logic_vector(31 downto 0);
    signal conv80_2513 : std_logic_vector(31 downto 0);
    signal div5_2426 : std_logic_vector(15 downto 0);
    signal div98_2721 : std_logic_vector(15 downto 0);
    signal div_2408 : std_logic_vector(15 downto 0);
    signal iNsTr_10_2505 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2398 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2416 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2434 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2444 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2456 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2469 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2481 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2493 : std_logic_vector(31 downto 0);
    signal inc95_2715 : std_logic_vector(15 downto 0);
    signal inc_2704 : std_logic_vector(15 downto 0);
    signal indvar_2603 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2696 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2733 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2544 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2538 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2727 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2616 : std_logic_vector(15 downto 0);
    signal ptr_deref_2401_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2401_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2401_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2401_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2401_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2419_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2419_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2419_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2419_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2419_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2437_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2437_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2437_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2437_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2437_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2447_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2447_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2447_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2447_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2447_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2459_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2459_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2459_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2459_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2459_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2472_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2472_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2472_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2472_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2472_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2484_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2484_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2484_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2484_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2484_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2496_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2496_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2496_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2496_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2496_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2508_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2508_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2508_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2508_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2508_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2646_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2646_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2646_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2646_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2646_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2666_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2666_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2666_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2666_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2666_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2666_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr118_2636 : std_logic_vector(63 downto 0);
    signal shr72120_2657 : std_logic_vector(63 downto 0);
    signal tmp10_2580 : std_logic_vector(15 downto 0);
    signal tmp11_2585 : std_logic_vector(15 downto 0);
    signal tmp12_2590 : std_logic_vector(15 downto 0);
    signal tmp134_2555 : std_logic_vector(15 downto 0);
    signal tmp135_2560 : std_logic_vector(15 downto 0);
    signal tmp136_2565 : std_logic_vector(15 downto 0);
    signal tmp13_2595 : std_logic_vector(15 downto 0);
    signal tmp14_2600 : std_logic_vector(15 downto 0);
    signal tmp16_2438 : std_logic_vector(15 downto 0);
    signal tmp29_2448 : std_logic_vector(15 downto 0);
    signal tmp32_2460 : std_logic_vector(15 downto 0);
    signal tmp35_2463 : std_logic_vector(15 downto 0);
    signal tmp3_2420 : std_logic_vector(15 downto 0);
    signal tmp41_2473 : std_logic_vector(15 downto 0);
    signal tmp44_2485 : std_logic_vector(15 downto 0);
    signal tmp4_2519 : std_logic_vector(15 downto 0);
    signal tmp54_2497 : std_logic_vector(15 downto 0);
    signal tmp58_2509 : std_logic_vector(15 downto 0);
    signal tmp5_2524 : std_logic_vector(15 downto 0);
    signal tmp69_2647 : std_logic_vector(63 downto 0);
    signal tmp6_2570 : std_logic_vector(15 downto 0);
    signal tmp7_2575 : std_logic_vector(15 downto 0);
    signal tmp8_2530 : std_logic_vector(15 downto 0);
    signal tmp9_2535 : std_logic_vector(15 downto 0);
    signal tmp_2402 : std_logic_vector(15 downto 0);
    signal type_cast_2406_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2424_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2517_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2528_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2541_wire : std_logic_vector(15 downto 0);
    signal type_cast_2543_wire : std_logic_vector(15 downto 0);
    signal type_cast_2547_wire : std_logic_vector(15 downto 0);
    signal type_cast_2549_wire : std_logic_vector(15 downto 0);
    signal type_cast_2607_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2609_wire : std_logic_vector(15 downto 0);
    signal type_cast_2614_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2634_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2655_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2676_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2694_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2702_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2713_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2719_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    LOAD_padding_2462_word_address_0 <= "0";
    array_obj_ref_2641_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2641_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2641_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2641_resized_base_address <= "00000000000000";
    array_obj_ref_2662_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2662_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2662_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2662_resized_base_address <= "00000000000000";
    iNsTr_10_2505 <= "00000000000000000000000000000100";
    iNsTr_2_2398 <= "00000000000000000000000000000011";
    iNsTr_3_2416 <= "00000000000000000000000000000100";
    iNsTr_4_2434 <= "00000000000000000000000000000101";
    iNsTr_5_2444 <= "00000000000000000000000000000000";
    iNsTr_6_2456 <= "00000000000000000000000000000100";
    iNsTr_7_2469 <= "00000000000000000000000000000001";
    iNsTr_8_2481 <= "00000000000000000000000000000101";
    iNsTr_9_2493 <= "00000000000000000000000000000101";
    ptr_deref_2401_word_offset_0 <= "0000000";
    ptr_deref_2419_word_offset_0 <= "0000000";
    ptr_deref_2437_word_offset_0 <= "0000000";
    ptr_deref_2447_word_offset_0 <= "0";
    ptr_deref_2459_word_offset_0 <= "0000000";
    ptr_deref_2472_word_offset_0 <= "0";
    ptr_deref_2484_word_offset_0 <= "0000000";
    ptr_deref_2496_word_offset_0 <= "0000000";
    ptr_deref_2508_word_offset_0 <= "0000000";
    ptr_deref_2646_word_offset_0 <= "00000000000000";
    ptr_deref_2666_word_offset_0 <= "00000000000000";
    type_cast_2406_wire_constant <= "0000000000000001";
    type_cast_2424_wire_constant <= "0000000000000001";
    type_cast_2517_wire_constant <= "1111111111111111";
    type_cast_2528_wire_constant <= "1111111111111111";
    type_cast_2607_wire_constant <= "0000000000000000";
    type_cast_2614_wire_constant <= "0000000000000100";
    type_cast_2634_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2655_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2676_wire_constant <= "00000000000000000000000000000100";
    type_cast_2694_wire_constant <= "0000000000000001";
    type_cast_2702_wire_constant <= "0000000000000001";
    type_cast_2713_wire_constant <= "0000000000000001";
    type_cast_2719_wire_constant <= "0000000000000001";
    phi_stmt_2538: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2541_wire & type_cast_2543_wire;
      req <= phi_stmt_2538_req_0 & phi_stmt_2538_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2538",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2538_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2538,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2538
    phi_stmt_2544: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2547_wire & type_cast_2549_wire;
      req <= phi_stmt_2544_req_0 & phi_stmt_2544_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2544",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2544_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2544,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2544
    phi_stmt_2603: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2607_wire_constant & type_cast_2609_wire;
      req <= phi_stmt_2603_req_0 & phi_stmt_2603_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2603",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2603_ack_0,
          idata => idata,
          odata => indvar_2603,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2603
    -- flow-through select operator MUX_2726_inst
    input_dim1x_x2_2727 <= div98_2721 when (cmp91_2709(0) /=  '0') else inc_2704;
    -- flow-through select operator MUX_2732_inst
    input_dim0x_x0_2733 <= inc95_2715 when (cmp91_2709(0) /=  '0') else input_dim0x_x2x_xph_2544;
    addr_of_2642_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2642_final_reg_req_0;
      addr_of_2642_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2642_final_reg_req_1;
      addr_of_2642_final_reg_ack_1<= rack(0);
      addr_of_2642_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2642_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2641_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2643,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2663_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2663_final_reg_req_0;
      addr_of_2663_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2663_final_reg_req_1;
      addr_of_2663_final_reg_ack_1<= rack(0);
      addr_of_2663_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2663_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2662_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx74_2664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2512_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2512_inst_req_0;
      type_cast_2512_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2512_inst_req_1;
      type_cast_2512_inst_ack_1<= rack(0);
      type_cast_2512_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2512_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp16_2438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2513,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2541_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2541_inst_req_0;
      type_cast_2541_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2541_inst_req_1;
      type_cast_2541_inst_ack_1<= rack(0);
      type_cast_2541_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2541_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2727,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2541_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2543_inst_req_0;
      type_cast_2543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2543_inst_req_1;
      type_cast_2543_inst_ack_1<= rack(0);
      type_cast_2543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div5_2426,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2543_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2547_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2547_inst_req_0;
      type_cast_2547_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2547_inst_req_1;
      type_cast_2547_inst_ack_1<= rack(0);
      type_cast_2547_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2547_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2408,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2547_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2549_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2549_inst_req_0;
      type_cast_2549_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2549_inst_req_1;
      type_cast_2549_inst_ack_1<= rack(0);
      type_cast_2549_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2549_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2733,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2549_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2609_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2609_inst_req_0;
      type_cast_2609_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2609_inst_req_1;
      type_cast_2609_inst_ack_1<= rack(0);
      type_cast_2609_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2609_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2696,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2609_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2629_inst_req_0;
      type_cast_2629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2629_inst_req_1;
      type_cast_2629_inst_ack_1<= rack(0);
      type_cast_2629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2629_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add25_2621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2630,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2650_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2650_inst_req_0;
      type_cast_2650_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2650_inst_req_1;
      type_cast_2650_inst_ack_1<= rack(0);
      type_cast_2650_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2650_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add65_2626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_2651,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2671_inst_req_0;
      type_cast_2671_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2671_inst_req_1;
      type_cast_2671_inst_ack_1<= rack(0);
      type_cast_2671_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2671_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2616,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv77_2672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2462_gather_scatter
    process(LOAD_padding_2462_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2462_data_0;
      ov(15 downto 0) := iv;
      tmp35_2463 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2641_index_1_rename
    process(R_shr118_2640_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr118_2640_resized;
      ov(13 downto 0) := iv;
      R_shr118_2640_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2641_index_1_resize
    process(shr118_2636) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr118_2636;
      ov := iv(13 downto 0);
      R_shr118_2640_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2641_root_address_inst
    process(array_obj_ref_2641_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2641_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2641_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2662_index_1_rename
    process(R_shr72120_2661_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_shr72120_2661_resized;
      ov(13 downto 0) := iv;
      R_shr72120_2661_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2662_index_1_resize
    process(shr72120_2657) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shr72120_2657;
      ov := iv(13 downto 0);
      R_shr72120_2661_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2662_root_address_inst
    process(array_obj_ref_2662_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2662_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2662_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2401_addr_0
    process(ptr_deref_2401_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2401_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2401_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2401_base_resize
    process(iNsTr_2_2398) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2398;
      ov := iv(6 downto 0);
      ptr_deref_2401_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2401_gather_scatter
    process(ptr_deref_2401_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2401_data_0;
      ov(15 downto 0) := iv;
      tmp_2402 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2401_root_address_inst
    process(ptr_deref_2401_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2401_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2401_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2419_addr_0
    process(ptr_deref_2419_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2419_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2419_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2419_base_resize
    process(iNsTr_3_2416) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2416;
      ov := iv(6 downto 0);
      ptr_deref_2419_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2419_gather_scatter
    process(ptr_deref_2419_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2419_data_0;
      ov(15 downto 0) := iv;
      tmp3_2420 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2419_root_address_inst
    process(ptr_deref_2419_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2419_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2419_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2437_addr_0
    process(ptr_deref_2437_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2437_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2437_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2437_base_resize
    process(iNsTr_4_2434) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2434;
      ov := iv(6 downto 0);
      ptr_deref_2437_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2437_gather_scatter
    process(ptr_deref_2437_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2437_data_0;
      ov(15 downto 0) := iv;
      tmp16_2438 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2437_root_address_inst
    process(ptr_deref_2437_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2437_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2437_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2447_addr_0
    process(ptr_deref_2447_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2447_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2447_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2447_base_resize
    process(iNsTr_5_2444) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2444;
      ov := iv(0 downto 0);
      ptr_deref_2447_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2447_gather_scatter
    process(ptr_deref_2447_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2447_data_0;
      ov(15 downto 0) := iv;
      tmp29_2448 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2447_root_address_inst
    process(ptr_deref_2447_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2447_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2447_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2459_addr_0
    process(ptr_deref_2459_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2459_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2459_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2459_base_resize
    process(iNsTr_6_2456) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2456;
      ov := iv(6 downto 0);
      ptr_deref_2459_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2459_gather_scatter
    process(ptr_deref_2459_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2459_data_0;
      ov(15 downto 0) := iv;
      tmp32_2460 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2459_root_address_inst
    process(ptr_deref_2459_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2459_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2459_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2472_addr_0
    process(ptr_deref_2472_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2472_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2472_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2472_base_resize
    process(iNsTr_7_2469) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2469;
      ov := iv(0 downto 0);
      ptr_deref_2472_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2472_gather_scatter
    process(ptr_deref_2472_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2472_data_0;
      ov(15 downto 0) := iv;
      tmp41_2473 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2472_root_address_inst
    process(ptr_deref_2472_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2472_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2472_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2484_addr_0
    process(ptr_deref_2484_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2484_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2484_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2484_base_resize
    process(iNsTr_8_2481) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2481;
      ov := iv(6 downto 0);
      ptr_deref_2484_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2484_gather_scatter
    process(ptr_deref_2484_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2484_data_0;
      ov(15 downto 0) := iv;
      tmp44_2485 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2484_root_address_inst
    process(ptr_deref_2484_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2484_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2484_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2496_addr_0
    process(ptr_deref_2496_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2496_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2496_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2496_base_resize
    process(iNsTr_9_2493) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2493;
      ov := iv(6 downto 0);
      ptr_deref_2496_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2496_gather_scatter
    process(ptr_deref_2496_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2496_data_0;
      ov(15 downto 0) := iv;
      tmp54_2497 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2496_root_address_inst
    process(ptr_deref_2496_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2496_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2496_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2508_addr_0
    process(ptr_deref_2508_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2508_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2508_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2508_base_resize
    process(iNsTr_10_2505) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2505;
      ov := iv(6 downto 0);
      ptr_deref_2508_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2508_gather_scatter
    process(ptr_deref_2508_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2508_data_0;
      ov(15 downto 0) := iv;
      tmp58_2509 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2508_root_address_inst
    process(ptr_deref_2508_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2508_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2508_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2646_addr_0
    process(ptr_deref_2646_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2646_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2646_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2646_base_resize
    process(arrayidx_2643) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2643;
      ov := iv(13 downto 0);
      ptr_deref_2646_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2646_gather_scatter
    process(ptr_deref_2646_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2646_data_0;
      ov(63 downto 0) := iv;
      tmp69_2647 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2646_root_address_inst
    process(ptr_deref_2646_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2646_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2646_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2666_addr_0
    process(ptr_deref_2666_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2666_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2666_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2666_base_resize
    process(arrayidx74_2664) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx74_2664;
      ov := iv(13 downto 0);
      ptr_deref_2666_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2666_gather_scatter
    process(tmp69_2647) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp69_2647;
      ov(63 downto 0) := iv;
      ptr_deref_2666_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2666_root_address_inst
    process(ptr_deref_2666_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2666_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2666_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2684_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2683;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2684_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2684_branch_req_0,
          ack0 => if_stmt_2684_branch_ack_0,
          ack1 => if_stmt_2684_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2739_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp104_2738;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2739_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2739_branch_req_0,
          ack0 => if_stmt_2739_branch_ack_0,
          ack1 => if_stmt_2739_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2518_inst
    process(tmp44_2485) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp44_2485, type_cast_2517_wire_constant, tmp_var);
      tmp4_2519 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2529_inst
    process(tmp32_2460) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp32_2460, type_cast_2528_wire_constant, tmp_var);
      tmp8_2530 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2559_inst
    process(input_dim1x_x1x_xph_2538, tmp134_2555) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2538, tmp134_2555, tmp_var);
      tmp135_2560 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2574_inst
    process(tmp5_2524, tmp6_2570) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp5_2524, tmp6_2570, tmp_var);
      tmp7_2575 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2584_inst
    process(tmp9_2535, tmp10_2580) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_2535, tmp10_2580, tmp_var);
      tmp11_2585 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2594_inst
    process(tmp7_2575, tmp12_2590) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp7_2575, tmp12_2590, tmp_var);
      tmp13_2595 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2620_inst
    process(tmp136_2565, input_dim2x_x1_2616) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp136_2565, input_dim2x_x1_2616, tmp_var);
      add25_2621 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2625_inst
    process(tmp14_2600, input_dim2x_x1_2616) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp14_2600, input_dim2x_x1_2616, tmp_var);
      add65_2626 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2695_inst
    process(indvar_2603) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2603, type_cast_2694_wire_constant, tmp_var);
      indvarx_xnext_2696 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2703_inst
    process(input_dim1x_x1x_xph_2538) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2538, type_cast_2702_wire_constant, tmp_var);
      inc_2704 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2714_inst
    process(input_dim0x_x2x_xph_2544) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_2544, type_cast_2713_wire_constant, tmp_var);
      inc95_2715 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2677_inst
    process(conv77_2672) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv77_2672, type_cast_2676_wire_constant, tmp_var);
      add78_2678 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2708_inst
    process(inc_2704, tmp3_2420) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2704, tmp3_2420, tmp_var);
      cmp91_2709 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2737_inst
    process(input_dim0x_x0_2733, tmp_2402) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(input_dim0x_x0_2733, tmp_2402, tmp_var);
      cmp104_2738 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2407_inst
    process(tmp_2402) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2402, type_cast_2406_wire_constant, tmp_var);
      div_2408 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2425_inst
    process(tmp3_2420) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_2420, type_cast_2424_wire_constant, tmp_var);
      div5_2426 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2720_inst
    process(tmp3_2420) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_2420, type_cast_2719_wire_constant, tmp_var);
      div98_2721 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2635_inst
    process(conv68_2630) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv68_2630, type_cast_2634_wire_constant, tmp_var);
      shr118_2636 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2656_inst
    process(conv71_2651) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv71_2651, type_cast_2655_wire_constant, tmp_var);
      shr72120_2657 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2554_inst
    process(tmp3_2420, input_dim0x_x2x_xph_2544) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp3_2420, input_dim0x_x2x_xph_2544, tmp_var);
      tmp134_2555 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2564_inst
    process(tmp16_2438, tmp135_2560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_2438, tmp135_2560, tmp_var);
      tmp136_2565 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2569_inst
    process(tmp41_2473, input_dim1x_x1x_xph_2538) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp41_2473, input_dim1x_x1x_xph_2538, tmp_var);
      tmp6_2570 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2579_inst
    process(tmp29_2448, input_dim0x_x2x_xph_2544) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp29_2448, input_dim0x_x2x_xph_2544, tmp_var);
      tmp10_2580 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2589_inst
    process(tmp58_2509, tmp11_2585) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp58_2509, tmp11_2585, tmp_var);
      tmp12_2590 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2599_inst
    process(tmp54_2497, tmp13_2595) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_2497, tmp13_2595, tmp_var);
      tmp14_2600 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2615_inst
    process(indvar_2603) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2603, type_cast_2614_wire_constant, tmp_var);
      input_dim2x_x1_2616 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2523_inst
    process(tmp4_2519, tmp35_2463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp4_2519, tmp35_2463, tmp_var);
      tmp5_2524 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2534_inst
    process(tmp8_2530, tmp35_2463) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(tmp8_2530, tmp35_2463, tmp_var);
      tmp9_2535 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2682_inst
    process(add78_2678, conv80_2513) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add78_2678, conv80_2513, tmp_var);
      cmp_2683 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2641_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr118_2640_scaled;
      array_obj_ref_2641_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2641_index_offset_req_0;
      array_obj_ref_2641_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2641_index_offset_req_1;
      array_obj_ref_2641_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2662_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_shr72120_2661_scaled;
      array_obj_ref_2662_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2662_index_offset_req_0;
      array_obj_ref_2662_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2662_index_offset_req_1;
      array_obj_ref_2662_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : LOAD_padding_2462_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2462_load_0_req_0;
      LOAD_padding_2462_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2462_load_0_req_1;
      LOAD_padding_2462_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2462_word_address_0;
      LOAD_padding_2462_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2401_load_0 ptr_deref_2437_load_0 ptr_deref_2419_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2401_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2437_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2419_load_0_req_0;
      ptr_deref_2401_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2437_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2419_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2401_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2437_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2419_load_0_req_1;
      ptr_deref_2401_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2437_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2419_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2401_word_address_0 & ptr_deref_2437_word_address_0 & ptr_deref_2419_word_address_0;
      ptr_deref_2401_data_0 <= data_out(47 downto 32);
      ptr_deref_2437_data_0 <= data_out(31 downto 16);
      ptr_deref_2419_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2447_load_0 ptr_deref_2472_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2447_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2472_load_0_req_0;
      ptr_deref_2447_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2472_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2447_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2472_load_0_req_1;
      ptr_deref_2447_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2472_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2447_word_address_0 & ptr_deref_2472_word_address_0;
      ptr_deref_2447_data_0 <= data_out(31 downto 16);
      ptr_deref_2472_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2459_load_0 ptr_deref_2484_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2459_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2484_load_0_req_0;
      ptr_deref_2459_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2484_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2459_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2484_load_0_req_1;
      ptr_deref_2459_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2484_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2459_word_address_0 & ptr_deref_2484_word_address_0;
      ptr_deref_2459_data_0 <= data_out(31 downto 16);
      ptr_deref_2484_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2508_load_0 ptr_deref_2496_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2508_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2496_load_0_req_0;
      ptr_deref_2508_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2496_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2508_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2496_load_0_req_1;
      ptr_deref_2508_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2496_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2508_word_address_0 & ptr_deref_2496_word_address_0;
      ptr_deref_2508_data_0 <= data_out(31 downto 16);
      ptr_deref_2496_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2646_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2646_load_0_req_0;
      ptr_deref_2646_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2646_load_0_req_1;
      ptr_deref_2646_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2646_word_address_0;
      ptr_deref_2646_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2666_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2666_store_0_req_0;
      ptr_deref_2666_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2666_store_0_req_1;
      ptr_deref_2666_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2666_word_address_0;
      data_in <= ptr_deref_2666_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2388_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_start_2388_inst_req_0;
      RPIPE_Block3_start_2388_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_start_2388_inst_req_1;
      RPIPE_Block3_start_2388_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2389 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2747_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2747_inst_req_0;
      WPIPE_Block3_done_2747_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2747_inst_req_1;
      WPIPE_Block3_done_2747_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2389;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_2934_start: Boolean;
  signal sendOutput_CP_2934_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_984_load_0_req_1 : boolean;
  signal ptr_deref_984_load_0_ack_1 : boolean;
  signal type_cast_988_inst_req_0 : boolean;
  signal type_cast_988_inst_ack_0 : boolean;
  signal ptr_deref_984_load_0_req_0 : boolean;
  signal ptr_deref_984_load_0_ack_0 : boolean;
  signal type_cast_988_inst_req_1 : boolean;
  signal type_cast_988_inst_ack_1 : boolean;
  signal type_cast_1004_inst_req_0 : boolean;
  signal type_cast_1004_inst_ack_0 : boolean;
  signal type_cast_1004_inst_req_1 : boolean;
  signal type_cast_1004_inst_ack_1 : boolean;
  signal ptr_deref_1000_load_0_req_1 : boolean;
  signal ptr_deref_1000_load_0_ack_1 : boolean;
  signal ptr_deref_1000_load_0_req_0 : boolean;
  signal ptr_deref_1000_load_0_ack_0 : boolean;
  signal phi_stmt_1081_ack_0 : boolean;
  signal ptr_deref_1016_load_0_req_0 : boolean;
  signal ptr_deref_1016_load_0_ack_0 : boolean;
  signal ptr_deref_1016_load_0_req_1 : boolean;
  signal ptr_deref_1016_load_0_ack_1 : boolean;
  signal type_cast_1020_inst_req_0 : boolean;
  signal type_cast_1020_inst_ack_0 : boolean;
  signal type_cast_1020_inst_req_1 : boolean;
  signal type_cast_1020_inst_ack_1 : boolean;
  signal if_stmt_1053_branch_req_0 : boolean;
  signal if_stmt_1053_branch_ack_1 : boolean;
  signal if_stmt_1053_branch_ack_0 : boolean;
  signal array_obj_ref_1093_index_offset_req_0 : boolean;
  signal array_obj_ref_1093_index_offset_ack_0 : boolean;
  signal array_obj_ref_1093_index_offset_req_1 : boolean;
  signal array_obj_ref_1093_index_offset_ack_1 : boolean;
  signal addr_of_1094_final_reg_req_0 : boolean;
  signal addr_of_1094_final_reg_ack_0 : boolean;
  signal addr_of_1094_final_reg_req_1 : boolean;
  signal addr_of_1094_final_reg_ack_1 : boolean;
  signal ptr_deref_1098_load_0_req_0 : boolean;
  signal ptr_deref_1098_load_0_ack_0 : boolean;
  signal ptr_deref_1098_load_0_req_1 : boolean;
  signal ptr_deref_1098_load_0_ack_1 : boolean;
  signal type_cast_1102_inst_req_0 : boolean;
  signal type_cast_1102_inst_ack_0 : boolean;
  signal type_cast_1102_inst_req_1 : boolean;
  signal type_cast_1102_inst_ack_1 : boolean;
  signal type_cast_1112_inst_req_0 : boolean;
  signal type_cast_1112_inst_ack_0 : boolean;
  signal type_cast_1112_inst_req_1 : boolean;
  signal type_cast_1112_inst_ack_1 : boolean;
  signal type_cast_1122_inst_req_0 : boolean;
  signal type_cast_1122_inst_ack_0 : boolean;
  signal type_cast_1122_inst_req_1 : boolean;
  signal type_cast_1122_inst_ack_1 : boolean;
  signal type_cast_1132_inst_req_0 : boolean;
  signal type_cast_1132_inst_ack_0 : boolean;
  signal type_cast_1132_inst_req_1 : boolean;
  signal type_cast_1132_inst_ack_1 : boolean;
  signal type_cast_1142_inst_req_0 : boolean;
  signal type_cast_1142_inst_ack_0 : boolean;
  signal type_cast_1142_inst_req_1 : boolean;
  signal type_cast_1142_inst_ack_1 : boolean;
  signal type_cast_1152_inst_req_0 : boolean;
  signal type_cast_1152_inst_ack_0 : boolean;
  signal type_cast_1152_inst_req_1 : boolean;
  signal type_cast_1152_inst_ack_1 : boolean;
  signal type_cast_1162_inst_req_0 : boolean;
  signal type_cast_1162_inst_ack_0 : boolean;
  signal type_cast_1162_inst_req_1 : boolean;
  signal type_cast_1162_inst_ack_1 : boolean;
  signal type_cast_1172_inst_req_0 : boolean;
  signal type_cast_1172_inst_ack_0 : boolean;
  signal type_cast_1172_inst_req_1 : boolean;
  signal type_cast_1172_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1174_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1174_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1174_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1174_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1177_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1177_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1177_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1177_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1180_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1180_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1180_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1180_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1183_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1183_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1183_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1183_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1186_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1186_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1186_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1186_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1189_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1189_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1189_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1189_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1192_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1192_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1192_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1192_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1195_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1195_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1195_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1195_inst_ack_1 : boolean;
  signal if_stmt_1209_branch_req_0 : boolean;
  signal if_stmt_1209_branch_ack_1 : boolean;
  signal if_stmt_1209_branch_ack_0 : boolean;
  signal phi_stmt_1081_req_0 : boolean;
  signal type_cast_1087_inst_req_0 : boolean;
  signal type_cast_1087_inst_ack_0 : boolean;
  signal type_cast_1087_inst_req_1 : boolean;
  signal type_cast_1087_inst_ack_1 : boolean;
  signal phi_stmt_1081_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_2934_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_2934_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_2934_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_2934_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_2934: Block -- control-path 
    signal sendOutput_CP_2934_elements: BooleanArray(70 downto 0);
    -- 
  begin -- 
    sendOutput_CP_2934_elements(0) <= sendOutput_CP_2934_start;
    sendOutput_CP_2934_symbol <= sendOutput_CP_2934_elements(70);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (92) 
      -- CP-element group 0: 	 branch_block_stmt_973/branch_block_stmt_973__entry__
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052__entry__
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_update_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_update_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_973/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_update_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_update_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_update_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_update_start_
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_Update/cr
      -- 
    cr_3008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => ptr_deref_984_load_0_req_1); -- 
    rr_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => ptr_deref_984_load_0_req_0); -- 
    cr_3027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => type_cast_988_inst_req_1); -- 
    cr_3091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => type_cast_1004_inst_req_1); -- 
    cr_3072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => ptr_deref_1000_load_0_req_1); -- 
    rr_3061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => ptr_deref_1000_load_0_req_0); -- 
    rr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => ptr_deref_1016_load_0_req_0); -- 
    cr_3136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => ptr_deref_1016_load_0_req_1); -- 
    cr_3155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(0), ack => type_cast_1020_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Sample/word_access_start/word_0/ra
      -- 
    ra_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_984_load_0_ack_0, ack => sendOutput_CP_2934_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (12) 
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/ptr_deref_984_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/ptr_deref_984_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/ptr_deref_984_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_984_Update/ptr_deref_984_Merge/merge_ack
      -- 
    ca_3009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_984_load_0_ack_1, ack => sendOutput_CP_2934_elements(2)); -- 
    rr_3022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(2), ack => type_cast_988_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_Sample/$exit
      -- 
    ra_3023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_988_inst_ack_0, ack => sendOutput_CP_2934_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	13 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_988_Update/ca
      -- 
    ca_3028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_988_inst_ack_1, ack => sendOutput_CP_2934_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Sample/word_access_start/word_0/ra
      -- 
    ra_3062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1000_load_0_ack_0, ack => sendOutput_CP_2934_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (12) 
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/ptr_deref_1000_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/ptr_deref_1000_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/ptr_deref_1000_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/ptr_deref_1000_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1000_Update/word_access_complete/$exit
      -- 
    ca_3073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1000_load_0_ack_1, ack => sendOutput_CP_2934_elements(6)); -- 
    rr_3086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(6), ack => type_cast_1004_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_Sample/ra
      -- 
    ra_3087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1004_inst_ack_0, ack => sendOutput_CP_2934_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1004_Update/ca
      -- 
    ca_3092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1004_inst_ack_1, ack => sendOutput_CP_2934_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Sample/word_access_start/word_0/ra
      -- 
    ra_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_0_ack_0, ack => sendOutput_CP_2934_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/ptr_deref_1016_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/ptr_deref_1016_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/ptr_deref_1016_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/ptr_deref_1016_Update/ptr_deref_1016_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_Sample/rr
      -- 
    ca_3137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1016_load_0_ack_1, ack => sendOutput_CP_2934_elements(10)); -- 
    rr_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(10), ack => type_cast_1020_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_Sample/ra
      -- 
    ra_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1020_inst_ack_0, ack => sendOutput_CP_2934_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/type_cast_1020_Update/ca
      -- 
    ca_3156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1020_inst_ack_1, ack => sendOutput_CP_2934_elements(12)); -- 
    -- CP-element group 13:  branch  join  transition  place  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: 	4 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (10) 
      -- CP-element group 13: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052/$exit
      -- CP-element group 13: 	 branch_block_stmt_973/assign_stmt_981_to_assign_stmt_1052__exit__
      -- CP-element group 13: 	 branch_block_stmt_973/if_stmt_1053__entry__
      -- CP-element group 13: 	 branch_block_stmt_973/if_stmt_1053_dead_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_973/if_stmt_1053_eval_test/$entry
      -- CP-element group 13: 	 branch_block_stmt_973/if_stmt_1053_eval_test/$exit
      -- CP-element group 13: 	 branch_block_stmt_973/if_stmt_1053_eval_test/branch_req
      -- CP-element group 13: 	 branch_block_stmt_973/R_cmp80_1054_place
      -- CP-element group 13: 	 branch_block_stmt_973/if_stmt_1053_if_link/$entry
      -- CP-element group 13: 	 branch_block_stmt_973/if_stmt_1053_else_link/$entry
      -- 
    branch_req_3164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(13), ack => if_stmt_1053_branch_req_0); -- 
    sendOutput_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(12) & sendOutput_CP_2934_elements(4) & sendOutput_CP_2934_elements(8);
      gj_sendOutput_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  merge  transition  place  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	64 
    -- CP-element group 14:  members (18) 
      -- CP-element group 14: 	 branch_block_stmt_973/bbx_xnph_forx_xbody
      -- CP-element group 14: 	 branch_block_stmt_973/assign_stmt_1065_to_assign_stmt_1078__exit__
      -- CP-element group 14: 	 branch_block_stmt_973/merge_stmt_1059__exit__
      -- CP-element group 14: 	 branch_block_stmt_973/assign_stmt_1065_to_assign_stmt_1078__entry__
      -- CP-element group 14: 	 branch_block_stmt_973/if_stmt_1053_if_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_973/if_stmt_1053_if_link/if_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_973/entry_bbx_xnph
      -- CP-element group 14: 	 branch_block_stmt_973/assign_stmt_1065_to_assign_stmt_1078/$entry
      -- CP-element group 14: 	 branch_block_stmt_973/assign_stmt_1065_to_assign_stmt_1078/$exit
      -- CP-element group 14: 	 branch_block_stmt_973/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_973/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_973/merge_stmt_1059_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_973/merge_stmt_1059_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_973/merge_stmt_1059_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_973/merge_stmt_1059_PhiAck/dummy
      -- CP-element group 14: 	 branch_block_stmt_973/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_973/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1081/$entry
      -- CP-element group 14: 	 branch_block_stmt_973/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/$entry
      -- 
    if_choice_transition_3169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1053_branch_ack_1, ack => sendOutput_CP_2934_elements(14)); -- 
    -- CP-element group 15:  transition  place  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	70 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_973/entry_forx_xend_PhiReq/$exit
      -- CP-element group 15: 	 branch_block_stmt_973/entry_forx_xend_PhiReq/$entry
      -- CP-element group 15: 	 branch_block_stmt_973/if_stmt_1053_else_link/$exit
      -- CP-element group 15: 	 branch_block_stmt_973/if_stmt_1053_else_link/else_choice_transition
      -- CP-element group 15: 	 branch_block_stmt_973/entry_forx_xend
      -- 
    else_choice_transition_3173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1053_branch_ack_0, ack => sendOutput_CP_2934_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	69 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	61 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_sample_complete
      -- CP-element group 16: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_Sample/ack
      -- 
    ack_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1093_index_offset_ack_0, ack => sendOutput_CP_2934_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	69 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (11) 
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_root_address_calculated
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_offset_calculated
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_Update/ack
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_base_plus_offset/$entry
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_base_plus_offset/$exit
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_base_plus_offset/sum_rename_req
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_base_plus_offset/sum_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_request/$entry
      -- CP-element group 17: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_request/req
      -- 
    ack_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1093_index_offset_ack_1, ack => sendOutput_CP_2934_elements(17)); -- 
    req_3221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(17), ack => addr_of_1094_final_reg_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_request/$exit
      -- CP-element group 18: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_request/ack
      -- 
    ack_3222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1094_final_reg_ack_0, ack => sendOutput_CP_2934_elements(18)); -- 
    -- CP-element group 19:  join  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	69 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (24) 
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_complete/$exit
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_complete/ack
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_word_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_root_address_calculated
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_address_resized
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_addr_resize/$entry
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_addr_resize/$exit
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_addr_resize/base_resize_req
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_addr_resize/base_resize_ack
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_plus_offset/$entry
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_plus_offset/$exit
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_base_plus_offset/sum_rename_ack
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_word_addrgen/$entry
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_word_addrgen/$exit
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_word_addrgen/root_register_req
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_word_addrgen/root_register_ack
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Sample/word_access_start/$entry
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Sample/word_access_start/word_0/$entry
      -- CP-element group 19: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Sample/word_access_start/word_0/rr
      -- 
    ack_3227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1094_final_reg_ack_1, ack => sendOutput_CP_2934_elements(19)); -- 
    rr_3260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(19), ack => ptr_deref_1098_load_0_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Sample/word_access_start/$exit
      -- CP-element group 20: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Sample/word_access_start/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Sample/word_access_start/word_0/ra
      -- 
    ra_3261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1098_load_0_ack_0, ack => sendOutput_CP_2934_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	69 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	28 
    -- CP-element group 21: 	30 
    -- CP-element group 21: 	32 
    -- CP-element group 21: 	34 
    -- CP-element group 21: 	36 
    -- CP-element group 21:  members (33) 
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/word_access_complete/$exit
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/word_access_complete/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/word_access_complete/word_0/ca
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/ptr_deref_1098_Merge/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/ptr_deref_1098_Merge/$exit
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/ptr_deref_1098_Merge/merge_req
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/ptr_deref_1098_Merge/merge_ack
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_Sample/rr
      -- 
    ca_3272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1098_load_0_ack_1, ack => sendOutput_CP_2934_elements(21)); -- 
    rr_3299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(21), ack => type_cast_1112_inst_req_0); -- 
    rr_3313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(21), ack => type_cast_1122_inst_req_0); -- 
    rr_3327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(21), ack => type_cast_1132_inst_req_0); -- 
    rr_3341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(21), ack => type_cast_1142_inst_req_0); -- 
    rr_3355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(21), ack => type_cast_1152_inst_req_0); -- 
    rr_3369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(21), ack => type_cast_1162_inst_req_0); -- 
    rr_3383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(21), ack => type_cast_1172_inst_req_0); -- 
    rr_3285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(21), ack => type_cast_1102_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_Sample/ra
      -- 
    ra_3286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_0, ack => sendOutput_CP_2934_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	69 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	58 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_Update/ca
      -- 
    ca_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_1, ack => sendOutput_CP_2934_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_Sample/ra
      -- 
    ra_3300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_0, ack => sendOutput_CP_2934_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	69 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	55 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_Update/ca
      -- 
    ca_3305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_1, ack => sendOutput_CP_2934_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	21 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_Sample/ra
      -- 
    ra_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1122_inst_ack_0, ack => sendOutput_CP_2934_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	69 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	52 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_Update/ca
      -- 
    ca_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1122_inst_ack_1, ack => sendOutput_CP_2934_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	21 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_Sample/ra
      -- 
    ra_3328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1132_inst_ack_0, ack => sendOutput_CP_2934_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	69 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	49 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_Update/ca
      -- 
    ca_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1132_inst_ack_1, ack => sendOutput_CP_2934_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	21 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_Sample/ra
      -- 
    ra_3342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1142_inst_ack_0, ack => sendOutput_CP_2934_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	69 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	46 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_Update/ca
      -- 
    ca_3347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1142_inst_ack_1, ack => sendOutput_CP_2934_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	21 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_Sample/ra
      -- 
    ra_3356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1152_inst_ack_0, ack => sendOutput_CP_2934_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	69 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	43 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_Update/ca
      -- 
    ca_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1152_inst_ack_1, ack => sendOutput_CP_2934_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	21 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_Sample/ra
      -- 
    ra_3370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_0, ack => sendOutput_CP_2934_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	69 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	40 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_Update/ca
      -- 
    ca_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_1, ack => sendOutput_CP_2934_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	21 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_Sample/ra
      -- 
    ra_3384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1172_inst_ack_0, ack => sendOutput_CP_2934_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	69 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_Sample/req
      -- 
    ca_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1172_inst_ack_1, ack => sendOutput_CP_2934_elements(37)); -- 
    req_3397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(37), ack => WPIPE_ConvTranspose_output_pipe_1174_inst_req_0); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_update_start_
      -- CP-element group 38: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_Update/req
      -- 
    ack_3398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1174_inst_ack_0, ack => sendOutput_CP_2934_elements(38)); -- 
    req_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(38), ack => WPIPE_ConvTranspose_output_pipe_1174_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1174_Update/ack
      -- 
    ack_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1174_inst_ack_1, ack => sendOutput_CP_2934_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	35 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_Sample/req
      -- 
    req_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(40), ack => WPIPE_ConvTranspose_output_pipe_1177_inst_req_0); -- 
    sendOutput_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(35) & sendOutput_CP_2934_elements(39);
      gj_sendOutput_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_update_start_
      -- CP-element group 41: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_Sample/ack
      -- CP-element group 41: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_Update/req
      -- 
    ack_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1177_inst_ack_0, ack => sendOutput_CP_2934_elements(41)); -- 
    req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(41), ack => WPIPE_ConvTranspose_output_pipe_1177_inst_req_1); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1177_Update/ack
      -- 
    ack_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1177_inst_ack_1, ack => sendOutput_CP_2934_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	33 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_Sample/req
      -- 
    req_3425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(43), ack => WPIPE_ConvTranspose_output_pipe_1180_inst_req_0); -- 
    sendOutput_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(33) & sendOutput_CP_2934_elements(42);
      gj_sendOutput_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_update_start_
      -- CP-element group 44: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_Sample/ack
      -- CP-element group 44: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_Update/req
      -- 
    ack_3426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1180_inst_ack_0, ack => sendOutput_CP_2934_elements(44)); -- 
    req_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(44), ack => WPIPE_ConvTranspose_output_pipe_1180_inst_req_1); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1180_Update/ack
      -- 
    ack_3431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1180_inst_ack_1, ack => sendOutput_CP_2934_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	31 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_Sample/req
      -- 
    req_3439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(46), ack => WPIPE_ConvTranspose_output_pipe_1183_inst_req_0); -- 
    sendOutput_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(31) & sendOutput_CP_2934_elements(45);
      gj_sendOutput_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_update_start_
      -- CP-element group 47: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_Sample/ack
      -- CP-element group 47: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_Update/req
      -- 
    ack_3440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1183_inst_ack_0, ack => sendOutput_CP_2934_elements(47)); -- 
    req_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(47), ack => WPIPE_ConvTranspose_output_pipe_1183_inst_req_1); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1183_Update/ack
      -- 
    ack_3445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1183_inst_ack_1, ack => sendOutput_CP_2934_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	29 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_Sample/req
      -- 
    req_3453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(49), ack => WPIPE_ConvTranspose_output_pipe_1186_inst_req_0); -- 
    sendOutput_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(29) & sendOutput_CP_2934_elements(48);
      gj_sendOutput_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (6) 
      -- CP-element group 50: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_update_start_
      -- CP-element group 50: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_Update/req
      -- 
    ack_3454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1186_inst_ack_0, ack => sendOutput_CP_2934_elements(50)); -- 
    req_3458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(50), ack => WPIPE_ConvTranspose_output_pipe_1186_inst_req_1); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1186_Update/ack
      -- 
    ack_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1186_inst_ack_1, ack => sendOutput_CP_2934_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	27 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_Sample/req
      -- 
    req_3467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(52), ack => WPIPE_ConvTranspose_output_pipe_1189_inst_req_0); -- 
    sendOutput_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(27) & sendOutput_CP_2934_elements(51);
      gj_sendOutput_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_update_start_
      -- CP-element group 53: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_Sample/ack
      -- CP-element group 53: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_Update/req
      -- 
    ack_3468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1189_inst_ack_0, ack => sendOutput_CP_2934_elements(53)); -- 
    req_3472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(53), ack => WPIPE_ConvTranspose_output_pipe_1189_inst_req_1); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1189_Update/ack
      -- 
    ack_3473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1189_inst_ack_1, ack => sendOutput_CP_2934_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: 	25 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_Sample/req
      -- 
    req_3481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(55), ack => WPIPE_ConvTranspose_output_pipe_1192_inst_req_0); -- 
    sendOutput_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(54) & sendOutput_CP_2934_elements(25);
      gj_sendOutput_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_update_start_
      -- CP-element group 56: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_Sample/ack
      -- CP-element group 56: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_Update/req
      -- 
    ack_3482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1192_inst_ack_0, ack => sendOutput_CP_2934_elements(56)); -- 
    req_3486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(56), ack => WPIPE_ConvTranspose_output_pipe_1192_inst_req_1); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1192_Update/ack
      -- 
    ack_3487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1192_inst_ack_1, ack => sendOutput_CP_2934_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	23 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_Sample/req
      -- 
    req_3495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(58), ack => WPIPE_ConvTranspose_output_pipe_1195_inst_req_0); -- 
    sendOutput_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(23) & sendOutput_CP_2934_elements(57);
      gj_sendOutput_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_update_start_
      -- CP-element group 59: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_Update/req
      -- 
    ack_3496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1195_inst_ack_0, ack => sendOutput_CP_2934_elements(59)); -- 
    req_3500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(59), ack => WPIPE_ConvTranspose_output_pipe_1195_inst_req_1); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/WPIPE_ConvTranspose_output_pipe_1195_Update/ack
      -- 
    ack_3501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1195_inst_ack_1, ack => sendOutput_CP_2934_elements(60)); -- 
    -- CP-element group 61:  branch  join  transition  place  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	16 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (10) 
      -- CP-element group 61: 	 branch_block_stmt_973/if_stmt_1209__entry__
      -- CP-element group 61: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208__exit__
      -- CP-element group 61: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/$exit
      -- CP-element group 61: 	 branch_block_stmt_973/if_stmt_1209_dead_link/$entry
      -- CP-element group 61: 	 branch_block_stmt_973/if_stmt_1209_eval_test/$entry
      -- CP-element group 61: 	 branch_block_stmt_973/if_stmt_1209_eval_test/$exit
      -- CP-element group 61: 	 branch_block_stmt_973/if_stmt_1209_eval_test/branch_req
      -- CP-element group 61: 	 branch_block_stmt_973/R_exitcond4_1210_place
      -- CP-element group 61: 	 branch_block_stmt_973/if_stmt_1209_if_link/$entry
      -- CP-element group 61: 	 branch_block_stmt_973/if_stmt_1209_else_link/$entry
      -- 
    branch_req_3509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(61), ack => if_stmt_1209_branch_req_0); -- 
    sendOutput_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(16) & sendOutput_CP_2934_elements(60);
      gj_sendOutput_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  merge  transition  place  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	70 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_973/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_973/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_973/merge_stmt_1215_PhiAck/dummy
      -- CP-element group 62: 	 branch_block_stmt_973/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_973/merge_stmt_1215_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_973/merge_stmt_1215__exit__
      -- CP-element group 62: 	 branch_block_stmt_973/forx_xendx_xloopexit_forx_xend
      -- CP-element group 62: 	 branch_block_stmt_973/merge_stmt_1215_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_973/merge_stmt_1215_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_973/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_973/if_stmt_1209_if_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_973/if_stmt_1209_if_link/if_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_973/forx_xbody_forx_xendx_xloopexit
      -- 
    if_choice_transition_3514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1209_branch_ack_1, ack => sendOutput_CP_2934_elements(62)); -- 
    -- CP-element group 63:  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (12) 
      -- CP-element group 63: 	 branch_block_stmt_973/if_stmt_1209_else_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_973/if_stmt_1209_else_link/else_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/$entry
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/$entry
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/$entry
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/$entry
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1209_branch_ack_0, ack => sendOutput_CP_2934_elements(63)); -- 
    rr_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(63), ack => type_cast_1087_inst_req_0); -- 
    cr_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(63), ack => type_cast_1087_inst_req_1); -- 
    -- CP-element group 64:  transition  output  delay-element  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	14 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	68 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_973/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_973/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1081/$exit
      -- CP-element group 64: 	 branch_block_stmt_973/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/$exit
      -- CP-element group 64: 	 branch_block_stmt_973/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1085_konst_delay_trans
      -- CP-element group 64: 	 branch_block_stmt_973/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_req
      -- 
    phi_stmt_1081_req_3543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1081_req_3543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(64), ack => phi_stmt_1081_req_0); -- 
    -- Element group sendOutput_CP_2934_elements(64) is a control-delay.
    cp_element_64_delay: control_delay_element  generic map(name => " 64_delay", delay_value => 1)  port map(req => sendOutput_CP_2934_elements(14), ack => sendOutput_CP_2934_elements(64), clk => clk, reset =>reset);
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/Sample/ra
      -- 
    ra_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1087_inst_ack_0, ack => sendOutput_CP_2934_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/Update/ca
      -- 
    ca_3568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1087_inst_ack_1, ack => sendOutput_CP_2934_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/$exit
      -- CP-element group 67: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/$exit
      -- CP-element group 67: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/$exit
      -- CP-element group 67: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_sources/type_cast_1087/SplitProtocol/$exit
      -- CP-element group 67: 	 branch_block_stmt_973/forx_xbody_forx_xbody_PhiReq/phi_stmt_1081/phi_stmt_1081_req
      -- 
    phi_stmt_1081_req_3569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1081_req_3569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(67), ack => phi_stmt_1081_req_1); -- 
    sendOutput_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_2934_elements(65) & sendOutput_CP_2934_elements(66);
      gj_sendOutput_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_2934_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  merge  transition  place  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	64 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_973/merge_stmt_1080_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_973/merge_stmt_1080_PhiReqMerge
      -- 
    sendOutput_CP_2934_elements(68) <= OrReduce(sendOutput_CP_2934_elements(64) & sendOutput_CP_2934_elements(67));
    -- CP-element group 69:  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	16 
    -- CP-element group 69: 	17 
    -- CP-element group 69: 	23 
    -- CP-element group 69: 	25 
    -- CP-element group 69: 	27 
    -- CP-element group 69: 	29 
    -- CP-element group 69: 	31 
    -- CP-element group 69: 	33 
    -- CP-element group 69: 	35 
    -- CP-element group 69: 	37 
    -- CP-element group 69: 	19 
    -- CP-element group 69: 	21 
    -- CP-element group 69:  members (53) 
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208__entry__
      -- CP-element group 69: 	 branch_block_stmt_973/merge_stmt_1080__exit__
      -- CP-element group 69: 	 branch_block_stmt_973/merge_stmt_1080_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_973/merge_stmt_1080_PhiAck/phi_stmt_1081_ack
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_resized_1
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_scaled_1
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_computed_1
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_resize_1/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_resize_1/$exit
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_resize_1/index_resize_req
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_resize_1/index_resize_ack
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_scale_1/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_scale_1/$exit
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_scale_1/scale_rename_req
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_index_scale_1/scale_rename_ack
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_update_start
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_Sample/req
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/array_obj_ref_1093_final_index_sum_regn_Update/req
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_complete/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/addr_of_1094_complete/req
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/word_access_complete/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/word_access_complete/word_0/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/ptr_deref_1098_Update/word_access_complete/word_0/cr
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1102_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1112_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1122_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1132_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1142_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1152_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1162_Update/cr
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_update_start_
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_973/assign_stmt_1095_to_assign_stmt_1208/type_cast_1172_Update/cr
      -- 
    phi_stmt_1081_ack_3574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1081_ack_0, ack => sendOutput_CP_2934_elements(69)); -- 
    req_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => array_obj_ref_1093_index_offset_req_0); -- 
    req_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => array_obj_ref_1093_index_offset_req_1); -- 
    req_3226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => addr_of_1094_final_reg_req_1); -- 
    cr_3271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => ptr_deref_1098_load_0_req_1); -- 
    cr_3290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => type_cast_1102_inst_req_1); -- 
    cr_3304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => type_cast_1112_inst_req_1); -- 
    cr_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => type_cast_1122_inst_req_1); -- 
    cr_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => type_cast_1132_inst_req_1); -- 
    cr_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => type_cast_1142_inst_req_1); -- 
    cr_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => type_cast_1152_inst_req_1); -- 
    cr_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => type_cast_1162_inst_req_1); -- 
    cr_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_2934_elements(69), ack => type_cast_1172_inst_req_1); -- 
    -- CP-element group 70:  merge  transition  place  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	15 
    -- CP-element group 70: 	62 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (16) 
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1217_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1219_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_973/return___PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1219__exit__
      -- CP-element group 70: 	 branch_block_stmt_973/branch_block_stmt_973__exit__
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1219_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1217_PhiAck/dummy
      -- CP-element group 70: 	 $exit
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1219_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1217__exit__
      -- CP-element group 70: 	 branch_block_stmt_973/return__
      -- CP-element group 70: 	 branch_block_stmt_973/$exit
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1217_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1219_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_973/return___PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_973/merge_stmt_1217_PhiReqMerge
      -- 
    sendOutput_CP_2934_elements(70) <= OrReduce(sendOutput_CP_2934_elements(15) & sendOutput_CP_2934_elements(62));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1044_wire : std_logic_vector(63 downto 0);
    signal R_indvar_1092_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1092_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1093_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1093_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1093_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1093_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1093_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1093_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1095 : std_logic_vector(31 downto 0);
    signal cmp80_1052 : std_logic_vector(0 downto 0);
    signal conv17_1103 : std_logic_vector(7 downto 0);
    signal conv23_1113 : std_logic_vector(7 downto 0);
    signal conv29_1123 : std_logic_vector(7 downto 0);
    signal conv2_1005 : std_logic_vector(63 downto 0);
    signal conv35_1133 : std_logic_vector(7 downto 0);
    signal conv41_1143 : std_logic_vector(7 downto 0);
    signal conv47_1153 : std_logic_vector(7 downto 0);
    signal conv4_1021 : std_logic_vector(63 downto 0);
    signal conv53_1163 : std_logic_vector(7 downto 0);
    signal conv59_1173 : std_logic_vector(7 downto 0);
    signal conv6_1046 : std_logic_vector(63 downto 0);
    signal conv_989 : std_logic_vector(63 downto 0);
    signal exitcond4_1208 : std_logic_vector(0 downto 0);
    signal iNsTr_0_981 : std_logic_vector(31 downto 0);
    signal iNsTr_1_997 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1013 : std_logic_vector(31 downto 0);
    signal indvar_1081 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1203 : std_logic_vector(63 downto 0);
    signal mul5_1032 : std_logic_vector(63 downto 0);
    signal mul_1027 : std_logic_vector(63 downto 0);
    signal ptr_deref_1000_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1000_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1000_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1000_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1000_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1016_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1016_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1016_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1016_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1016_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1098_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1098_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1098_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1098_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1098_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_984_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_984_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_984_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_984_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_984_word_offset_0 : std_logic_vector(6 downto 0);
    signal sext_1037 : std_logic_vector(63 downto 0);
    signal shr20_1109 : std_logic_vector(63 downto 0);
    signal shr26_1119 : std_logic_vector(63 downto 0);
    signal shr32_1129 : std_logic_vector(63 downto 0);
    signal shr38_1139 : std_logic_vector(63 downto 0);
    signal shr44_1149 : std_logic_vector(63 downto 0);
    signal shr50_1159 : std_logic_vector(63 downto 0);
    signal shr56_1169 : std_logic_vector(63 downto 0);
    signal shr_1065 : std_logic_vector(63 downto 0);
    signal tmp14_1099 : std_logic_vector(63 downto 0);
    signal tmp1_1001 : std_logic_vector(15 downto 0);
    signal tmp2_1071 : std_logic_vector(0 downto 0);
    signal tmp3_1017 : std_logic_vector(15 downto 0);
    signal tmp_985 : std_logic_vector(15 downto 0);
    signal type_cast_1025_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1040_wire : std_logic_vector(63 downto 0);
    signal type_cast_1043_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1050_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1063_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1069_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1076_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1085_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1087_wire : std_logic_vector(63 downto 0);
    signal type_cast_1107_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1117_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1127_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1137_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1147_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1157_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1167_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1201_wire_constant : std_logic_vector(63 downto 0);
    signal umax3_1078 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1093_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1093_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1093_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1093_resized_base_address <= "00000000000000";
    iNsTr_0_981 <= "00000000000000000000000000000011";
    iNsTr_1_997 <= "00000000000000000000000000000100";
    iNsTr_2_1013 <= "00000000000000000000000000000101";
    ptr_deref_1000_word_offset_0 <= "0000000";
    ptr_deref_1016_word_offset_0 <= "0000000";
    ptr_deref_1098_word_offset_0 <= "00000000000000";
    ptr_deref_984_word_offset_0 <= "0000000";
    type_cast_1025_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1043_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1050_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1063_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1069_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1076_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1085_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1107_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1117_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1127_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1137_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1147_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1157_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1167_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1201_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1081: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1085_wire_constant & type_cast_1087_wire;
      req <= phi_stmt_1081_req_0 & phi_stmt_1081_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1081",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1081_ack_0,
          idata => idata,
          odata => indvar_1081,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1081
    -- flow-through select operator MUX_1077_inst
    umax3_1078 <= shr_1065 when (tmp2_1071(0) /=  '0') else type_cast_1076_wire_constant;
    addr_of_1094_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1094_final_reg_req_0;
      addr_of_1094_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1094_final_reg_req_1;
      addr_of_1094_final_reg_ack_1<= rack(0);
      addr_of_1094_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1094_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1093_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1004_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1004_inst_req_0;
      type_cast_1004_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1004_inst_req_1;
      type_cast_1004_inst_ack_1<= rack(0);
      type_cast_1004_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1004_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_1001,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_1005,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1020_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1020_inst_req_0;
      type_cast_1020_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1020_inst_req_1;
      type_cast_1020_inst_ack_1<= rack(0);
      type_cast_1020_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1020_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_1017,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_1021,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1040_inst
    process(sext_1037) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1037(63 downto 0);
      type_cast_1040_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1045_inst
    process(ASHR_i64_i64_1044_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1044_wire(63 downto 0);
      conv6_1046 <= tmp_var; -- 
    end process;
    type_cast_1087_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1087_inst_req_0;
      type_cast_1087_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1087_inst_req_1;
      type_cast_1087_inst_ack_1<= rack(0);
      type_cast_1087_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1087_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1203,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1087_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1102_inst_req_0;
      type_cast_1102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1102_inst_req_1;
      type_cast_1102_inst_ack_1<= rack(0);
      type_cast_1102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_1099,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1112_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1112_inst_req_0;
      type_cast_1112_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1112_inst_req_1;
      type_cast_1112_inst_ack_1<= rack(0);
      type_cast_1112_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1112_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr20_1109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_1113,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1122_inst_req_0;
      type_cast_1122_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1122_inst_req_1;
      type_cast_1122_inst_ack_1<= rack(0);
      type_cast_1122_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1122_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr26_1119,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1123,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1132_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1132_inst_req_0;
      type_cast_1132_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1132_inst_req_1;
      type_cast_1132_inst_ack_1<= rack(0);
      type_cast_1132_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1132_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr32_1129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_1133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1142_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1142_inst_req_0;
      type_cast_1142_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1142_inst_req_1;
      type_cast_1142_inst_ack_1<= rack(0);
      type_cast_1142_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1142_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr38_1139,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_1143,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1152_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1152_inst_req_0;
      type_cast_1152_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1152_inst_req_1;
      type_cast_1152_inst_ack_1<= rack(0);
      type_cast_1152_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1152_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr44_1149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_1153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1162_inst_req_0;
      type_cast_1162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1162_inst_req_1;
      type_cast_1162_inst_ack_1<= rack(0);
      type_cast_1162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr50_1159,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1163,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1172_inst_req_0;
      type_cast_1172_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1172_inst_req_1;
      type_cast_1172_inst_ack_1<= rack(0);
      type_cast_1172_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1172_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr56_1169,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_1173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_988_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_988_inst_req_0;
      type_cast_988_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_988_inst_req_1;
      type_cast_988_inst_ack_1<= rack(0);
      type_cast_988_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_988_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_985,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_989,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1093_index_1_rename
    process(R_indvar_1092_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1092_resized;
      ov(13 downto 0) := iv;
      R_indvar_1092_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1093_index_1_resize
    process(indvar_1081) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1081;
      ov := iv(13 downto 0);
      R_indvar_1092_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1093_root_address_inst
    process(array_obj_ref_1093_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1093_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1093_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1000_addr_0
    process(ptr_deref_1000_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1000_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1000_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1000_base_resize
    process(iNsTr_1_997) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_997;
      ov := iv(6 downto 0);
      ptr_deref_1000_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1000_gather_scatter
    process(ptr_deref_1000_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1000_data_0;
      ov(15 downto 0) := iv;
      tmp1_1001 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1000_root_address_inst
    process(ptr_deref_1000_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1000_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1000_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1016_addr_0
    process(ptr_deref_1016_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1016_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1016_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1016_base_resize
    process(iNsTr_2_1013) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1013;
      ov := iv(6 downto 0);
      ptr_deref_1016_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1016_gather_scatter
    process(ptr_deref_1016_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1016_data_0;
      ov(15 downto 0) := iv;
      tmp3_1017 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1016_root_address_inst
    process(ptr_deref_1016_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1016_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1016_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1098_addr_0
    process(ptr_deref_1098_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1098_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1098_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1098_base_resize
    process(arrayidx_1095) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1095;
      ov := iv(13 downto 0);
      ptr_deref_1098_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1098_gather_scatter
    process(ptr_deref_1098_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1098_data_0;
      ov(63 downto 0) := iv;
      tmp14_1099 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1098_root_address_inst
    process(ptr_deref_1098_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1098_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1098_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_984_addr_0
    process(ptr_deref_984_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_984_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_984_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_984_base_resize
    process(iNsTr_0_981) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_981;
      ov := iv(6 downto 0);
      ptr_deref_984_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_984_gather_scatter
    process(ptr_deref_984_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_984_data_0;
      ov(15 downto 0) := iv;
      tmp_985 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_984_root_address_inst
    process(ptr_deref_984_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_984_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_984_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1053_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp80_1052;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1053_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1053_branch_req_0,
          ack0 => if_stmt_1053_branch_ack_0,
          ack1 => if_stmt_1053_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1209_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond4_1208;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1209_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1209_branch_req_0,
          ack0 => if_stmt_1209_branch_ack_0,
          ack1 => if_stmt_1209_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1202_inst
    process(indvar_1081) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1081, type_cast_1201_wire_constant, tmp_var);
      indvarx_xnext_1203 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1044_inst
    process(type_cast_1040_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1040_wire, type_cast_1043_wire_constant, tmp_var);
      ASHR_i64_i64_1044_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1207_inst
    process(indvarx_xnext_1203, umax3_1078) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1203, umax3_1078, tmp_var);
      exitcond4_1208 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1064_inst
    process(conv6_1046) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv6_1046, type_cast_1063_wire_constant, tmp_var);
      shr_1065 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1108_inst
    process(tmp14_1099) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_1099, type_cast_1107_wire_constant, tmp_var);
      shr20_1109 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1118_inst
    process(tmp14_1099) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_1099, type_cast_1117_wire_constant, tmp_var);
      shr26_1119 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1128_inst
    process(tmp14_1099) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_1099, type_cast_1127_wire_constant, tmp_var);
      shr32_1129 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1138_inst
    process(tmp14_1099) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_1099, type_cast_1137_wire_constant, tmp_var);
      shr38_1139 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1148_inst
    process(tmp14_1099) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_1099, type_cast_1147_wire_constant, tmp_var);
      shr44_1149 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1158_inst
    process(tmp14_1099) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_1099, type_cast_1157_wire_constant, tmp_var);
      shr50_1159 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1168_inst
    process(tmp14_1099) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_1099, type_cast_1167_wire_constant, tmp_var);
      shr56_1169 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1031_inst
    process(mul_1027, conv2_1005) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1027, conv2_1005, tmp_var);
      mul5_1032 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1036_inst
    process(mul5_1032, conv4_1021) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul5_1032, conv4_1021, tmp_var);
      sext_1037 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1026_inst
    process(conv_989) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_989, type_cast_1025_wire_constant, tmp_var);
      mul_1027 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1051_inst
    process(conv6_1046) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv6_1046, type_cast_1050_wire_constant, tmp_var);
      cmp80_1052 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1070_inst
    process(shr_1065) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_1065, type_cast_1069_wire_constant, tmp_var);
      tmp2_1071 <= tmp_var; --
    end process;
    -- shared split operator group (16) : array_obj_ref_1093_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1092_scaled;
      array_obj_ref_1093_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1093_index_offset_req_0;
      array_obj_ref_1093_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1093_index_offset_req_1;
      array_obj_ref_1093_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared load operator group (0) : ptr_deref_1016_load_0 ptr_deref_984_load_0 ptr_deref_1000_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1016_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_984_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1000_load_0_req_0;
      ptr_deref_1016_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_984_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1000_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1016_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_984_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1000_load_0_req_1;
      ptr_deref_1016_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_984_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1000_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1016_word_address_0 & ptr_deref_984_word_address_0 & ptr_deref_1000_word_address_0;
      ptr_deref_1016_data_0 <= data_out(47 downto 32);
      ptr_deref_984_data_0 <= data_out(31 downto 16);
      ptr_deref_1000_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(15 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1098_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1098_load_0_req_0;
      ptr_deref_1098_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1098_load_0_req_1;
      ptr_deref_1098_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1098_word_address_0;
      ptr_deref_1098_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(13 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(63 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1174_inst WPIPE_ConvTranspose_output_pipe_1186_inst WPIPE_ConvTranspose_output_pipe_1180_inst WPIPE_ConvTranspose_output_pipe_1183_inst WPIPE_ConvTranspose_output_pipe_1195_inst WPIPE_ConvTranspose_output_pipe_1177_inst WPIPE_ConvTranspose_output_pipe_1192_inst WPIPE_ConvTranspose_output_pipe_1189_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1174_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1186_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1180_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1183_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1195_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1177_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1192_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1189_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1174_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1186_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1180_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1183_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1195_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1177_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1192_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1189_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1174_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1186_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1180_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1183_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1195_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1177_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1192_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1189_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1174_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1186_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1180_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1183_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1195_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1177_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1192_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1189_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv59_1173 & conv35_1133 & conv47_1153 & conv41_1143 & conv17_1103 & conv53_1163 & conv23_1113 & conv29_1123;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_0_start: Boolean;
  signal testConfigure_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_933_inst_ack_1 : boolean;
  signal type_cast_861_inst_req_1 : boolean;
  signal ptr_deref_484_load_0_ack_1 : boolean;
  signal type_cast_504_inst_req_1 : boolean;
  signal type_cast_504_inst_ack_1 : boolean;
  signal type_cast_504_inst_req_0 : boolean;
  signal type_cast_160_inst_req_0 : boolean;
  signal type_cast_504_inst_ack_0 : boolean;
  signal phi_stmt_157_req_1 : boolean;
  signal type_cast_162_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_929_inst_req_0 : boolean;
  signal ptr_deref_381_store_0_ack_0 : boolean;
  signal type_cast_398_inst_ack_1 : boolean;
  signal ptr_deref_381_store_0_req_0 : boolean;
  signal type_cast_398_inst_req_1 : boolean;
  signal type_cast_398_inst_ack_0 : boolean;
  signal type_cast_398_inst_req_0 : boolean;
  signal type_cast_861_inst_ack_1 : boolean;
  signal ptr_deref_484_load_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal type_cast_472_inst_ack_1 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal type_cast_85_inst_req_0 : boolean;
  signal ptr_deref_394_load_0_ack_1 : boolean;
  signal ptr_deref_394_load_0_req_1 : boolean;
  signal ptr_deref_122_load_0_req_0 : boolean;
  signal ptr_deref_122_load_0_ack_0 : boolean;
  signal type_cast_370_inst_req_1 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_160_inst_req_1 : boolean;
  signal ptr_deref_47_store_0_req_0 : boolean;
  signal ptr_deref_47_store_0_ack_0 : boolean;
  signal ptr_deref_47_store_0_req_1 : boolean;
  signal ptr_deref_47_store_0_ack_1 : boolean;
  signal type_cast_915_inst_ack_1 : boolean;
  signal type_cast_370_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_req_1 : boolean;
  signal ptr_deref_426_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_929_inst_ack_0 : boolean;
  signal type_cast_62_inst_req_0 : boolean;
  signal ptr_deref_426_load_0_req_0 : boolean;
  signal type_cast_62_inst_ack_0 : boolean;
  signal type_cast_62_inst_req_1 : boolean;
  signal type_cast_62_inst_ack_1 : boolean;
  signal if_stmt_64_branch_req_0 : boolean;
  signal type_cast_472_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal if_stmt_64_branch_ack_1 : boolean;
  signal if_stmt_64_branch_ack_0 : boolean;
  signal type_cast_414_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_875_inst_req_0 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal ptr_deref_500_load_0_ack_1 : boolean;
  signal type_cast_488_inst_ack_1 : boolean;
  signal type_cast_414_inst_req_1 : boolean;
  signal array_obj_ref_101_index_offset_req_0 : boolean;
  signal array_obj_ref_101_index_offset_ack_0 : boolean;
  signal array_obj_ref_101_index_offset_req_1 : boolean;
  signal array_obj_ref_101_index_offset_ack_1 : boolean;
  signal ptr_deref_484_load_0_ack_0 : boolean;
  signal addr_of_102_final_reg_req_0 : boolean;
  signal addr_of_102_final_reg_ack_0 : boolean;
  signal addr_of_102_final_reg_req_1 : boolean;
  signal addr_of_102_final_reg_ack_1 : boolean;
  signal ptr_deref_500_load_0_req_1 : boolean;
  signal phi_stmt_157_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_875_inst_ack_0 : boolean;
  signal type_cast_430_inst_ack_1 : boolean;
  signal ptr_deref_484_load_0_req_0 : boolean;
  signal type_cast_160_inst_ack_1 : boolean;
  signal type_cast_488_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_929_inst_req_1 : boolean;
  signal ptr_deref_105_store_0_req_0 : boolean;
  signal ptr_deref_410_load_0_ack_1 : boolean;
  signal ptr_deref_105_store_0_ack_0 : boolean;
  signal ptr_deref_105_store_0_req_1 : boolean;
  signal ptr_deref_105_store_0_ack_1 : boolean;
  signal type_cast_430_inst_req_1 : boolean;
  signal type_cast_430_inst_ack_0 : boolean;
  signal type_cast_430_inst_req_0 : boolean;
  signal ptr_deref_410_load_0_req_1 : boolean;
  signal ptr_deref_381_store_0_ack_1 : boolean;
  signal ptr_deref_381_store_0_req_1 : boolean;
  signal addr_of_287_final_reg_req_0 : boolean;
  signal type_cast_897_inst_ack_0 : boolean;
  signal addr_of_287_final_reg_ack_0 : boolean;
  signal addr_of_287_final_reg_req_1 : boolean;
  signal addr_of_287_final_reg_ack_1 : boolean;
  signal type_cast_85_inst_ack_1 : boolean;
  signal phi_stmt_189_req_1 : boolean;
  signal ptr_deref_122_load_0_req_1 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal ptr_deref_122_load_0_ack_1 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_414_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal type_cast_915_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_137_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_137_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_137_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_137_inst_ack_1 : boolean;
  signal type_cast_141_inst_req_0 : boolean;
  signal type_cast_141_inst_ack_0 : boolean;
  signal type_cast_141_inst_req_1 : boolean;
  signal type_cast_141_inst_ack_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal if_stmt_143_branch_req_0 : boolean;
  signal if_stmt_143_branch_ack_1 : boolean;
  signal type_cast_414_inst_req_0 : boolean;
  signal if_stmt_143_branch_ack_0 : boolean;
  signal type_cast_85_inst_ack_0 : boolean;
  signal phi_stmt_73_req_0 : boolean;
  signal ptr_deref_171_store_0_req_0 : boolean;
  signal ptr_deref_171_store_0_ack_0 : boolean;
  signal ptr_deref_171_store_0_req_1 : boolean;
  signal ptr_deref_171_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_ack_1 : boolean;
  signal type_cast_370_inst_ack_0 : boolean;
  signal ptr_deref_468_load_0_ack_1 : boolean;
  signal if_stmt_180_branch_req_0 : boolean;
  signal type_cast_472_inst_ack_0 : boolean;
  signal ptr_deref_410_load_0_ack_0 : boolean;
  signal if_stmt_180_branch_ack_1 : boolean;
  signal if_stmt_180_branch_ack_0 : boolean;
  signal type_cast_205_inst_req_0 : boolean;
  signal type_cast_205_inst_ack_0 : boolean;
  signal ptr_deref_468_load_0_req_1 : boolean;
  signal type_cast_205_inst_req_1 : boolean;
  signal type_cast_205_inst_ack_1 : boolean;
  signal type_cast_472_inst_req_0 : boolean;
  signal type_cast_488_inst_ack_0 : boolean;
  signal ptr_deref_410_load_0_req_0 : boolean;
  signal type_cast_488_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_875_inst_ack_1 : boolean;
  signal array_obj_ref_211_index_offset_req_0 : boolean;
  signal array_obj_ref_211_index_offset_ack_0 : boolean;
  signal array_obj_ref_211_index_offset_req_1 : boolean;
  signal array_obj_ref_211_index_offset_ack_1 : boolean;
  signal addr_of_212_final_reg_req_0 : boolean;
  signal addr_of_212_final_reg_ack_0 : boolean;
  signal addr_of_212_final_reg_req_1 : boolean;
  signal addr_of_212_final_reg_ack_1 : boolean;
  signal ptr_deref_500_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_215_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_215_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_215_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_215_inst_ack_1 : boolean;
  signal type_cast_160_inst_ack_0 : boolean;
  signal type_cast_219_inst_req_0 : boolean;
  signal type_cast_219_inst_ack_0 : boolean;
  signal type_cast_219_inst_req_1 : boolean;
  signal type_cast_219_inst_ack_1 : boolean;
  signal ptr_deref_500_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_929_inst_ack_1 : boolean;
  signal type_cast_83_inst_req_1 : boolean;
  signal ptr_deref_394_load_0_ack_0 : boolean;
  signal phi_stmt_157_req_0 : boolean;
  signal ptr_deref_394_load_0_req_0 : boolean;
  signal ptr_deref_222_store_0_req_0 : boolean;
  signal ptr_deref_222_store_0_ack_0 : boolean;
  signal ptr_deref_222_store_0_req_1 : boolean;
  signal ptr_deref_222_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_875_inst_req_1 : boolean;
  signal ptr_deref_239_load_0_req_0 : boolean;
  signal ptr_deref_239_load_0_ack_0 : boolean;
  signal type_cast_370_inst_req_0 : boolean;
  signal ptr_deref_239_load_0_req_1 : boolean;
  signal ptr_deref_239_load_0_ack_1 : boolean;
  signal type_cast_243_inst_req_0 : boolean;
  signal type_cast_243_inst_ack_0 : boolean;
  signal type_cast_243_inst_req_1 : boolean;
  signal type_cast_243_inst_ack_1 : boolean;
  signal ptr_deref_468_load_0_ack_0 : boolean;
  signal if_stmt_252_branch_req_0 : boolean;
  signal type_cast_85_inst_req_1 : boolean;
  signal if_stmt_252_branch_ack_1 : boolean;
  signal if_stmt_252_branch_ack_0 : boolean;
  signal ptr_deref_468_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_ack_0 : boolean;
  signal ptr_deref_426_load_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_262_inst_ack_1 : boolean;
  signal type_cast_266_inst_req_0 : boolean;
  signal type_cast_266_inst_ack_0 : boolean;
  signal type_cast_266_inst_req_1 : boolean;
  signal type_cast_266_inst_ack_1 : boolean;
  signal ptr_deref_426_load_0_req_1 : boolean;
  signal phi_stmt_80_req_1 : boolean;
  signal ptr_deref_290_store_0_req_0 : boolean;
  signal ptr_deref_290_store_0_ack_0 : boolean;
  signal ptr_deref_290_store_0_req_1 : boolean;
  signal ptr_deref_290_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_294_inst_ack_1 : boolean;
  signal type_cast_298_inst_req_0 : boolean;
  signal type_cast_298_inst_ack_0 : boolean;
  signal type_cast_298_inst_req_1 : boolean;
  signal type_cast_298_inst_ack_1 : boolean;
  signal type_cast_897_inst_req_0 : boolean;
  signal if_stmt_312_branch_req_0 : boolean;
  signal if_stmt_312_branch_ack_1 : boolean;
  signal if_stmt_312_branch_ack_0 : boolean;
  signal STORE_padding_324_store_0_req_0 : boolean;
  signal STORE_padding_324_store_0_ack_0 : boolean;
  signal type_cast_83_inst_req_0 : boolean;
  signal STORE_padding_324_store_0_req_1 : boolean;
  signal type_cast_933_inst_req_0 : boolean;
  signal STORE_padding_324_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_ack_0 : boolean;
  signal type_cast_879_inst_req_0 : boolean;
  signal type_cast_83_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_328_inst_ack_1 : boolean;
  signal type_cast_879_inst_ack_0 : boolean;
  signal type_cast_332_inst_req_0 : boolean;
  signal type_cast_332_inst_ack_0 : boolean;
  signal type_cast_332_inst_req_1 : boolean;
  signal type_cast_332_inst_ack_1 : boolean;
  signal type_cast_933_inst_ack_0 : boolean;
  signal ptr_deref_343_store_0_req_0 : boolean;
  signal ptr_deref_343_store_0_ack_0 : boolean;
  signal ptr_deref_343_store_0_req_1 : boolean;
  signal ptr_deref_343_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_347_inst_ack_1 : boolean;
  signal type_cast_351_inst_req_0 : boolean;
  signal type_cast_351_inst_ack_0 : boolean;
  signal type_cast_351_inst_req_1 : boolean;
  signal type_cast_351_inst_ack_1 : boolean;
  signal ptr_deref_362_store_0_req_0 : boolean;
  signal ptr_deref_362_store_0_ack_0 : boolean;
  signal ptr_deref_362_store_0_req_1 : boolean;
  signal ptr_deref_362_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 : boolean;
  signal type_cast_966_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_893_inst_req_0 : boolean;
  signal ptr_deref_516_load_0_req_0 : boolean;
  signal type_cast_966_inst_req_1 : boolean;
  signal ptr_deref_516_load_0_ack_0 : boolean;
  signal type_cast_933_inst_req_1 : boolean;
  signal ptr_deref_516_load_0_req_1 : boolean;
  signal ptr_deref_516_load_0_ack_1 : boolean;
  signal type_cast_966_inst_ack_0 : boolean;
  signal type_cast_520_inst_req_0 : boolean;
  signal type_cast_520_inst_ack_0 : boolean;
  signal type_cast_520_inst_req_1 : boolean;
  signal type_cast_520_inst_ack_1 : boolean;
  signal type_cast_162_inst_req_1 : boolean;
  signal type_cast_966_inst_req_0 : boolean;
  signal phi_stmt_73_req_1 : boolean;
  signal if_stmt_558_branch_req_0 : boolean;
  signal if_stmt_558_branch_ack_1 : boolean;
  signal if_stmt_558_branch_ack_0 : boolean;
  signal phi_stmt_189_req_0 : boolean;
  signal if_stmt_573_branch_req_0 : boolean;
  signal if_stmt_573_branch_ack_1 : boolean;
  signal type_cast_879_inst_ack_1 : boolean;
  signal if_stmt_573_branch_ack_0 : boolean;
  signal type_cast_162_inst_ack_0 : boolean;
  signal type_cast_162_inst_req_0 : boolean;
  signal type_cast_879_inst_req_1 : boolean;
  signal phi_stmt_80_req_0 : boolean;
  signal type_cast_83_inst_ack_1 : boolean;
  signal array_obj_ref_613_index_offset_req_0 : boolean;
  signal array_obj_ref_613_index_offset_ack_0 : boolean;
  signal array_obj_ref_613_index_offset_req_1 : boolean;
  signal array_obj_ref_613_index_offset_ack_1 : boolean;
  signal if_stmt_955_branch_ack_0 : boolean;
  signal type_cast_915_inst_ack_0 : boolean;
  signal addr_of_614_final_reg_req_0 : boolean;
  signal addr_of_614_final_reg_ack_0 : boolean;
  signal addr_of_614_final_reg_req_1 : boolean;
  signal phi_stmt_150_ack_0 : boolean;
  signal addr_of_614_final_reg_ack_1 : boolean;
  signal type_cast_915_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_617_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_617_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_617_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_617_inst_ack_1 : boolean;
  signal type_cast_192_inst_ack_1 : boolean;
  signal type_cast_621_inst_req_0 : boolean;
  signal phi_stmt_150_req_0 : boolean;
  signal type_cast_621_inst_ack_0 : boolean;
  signal type_cast_621_inst_req_1 : boolean;
  signal type_cast_153_inst_ack_1 : boolean;
  signal type_cast_621_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_630_inst_req_0 : boolean;
  signal type_cast_153_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_630_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_630_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_630_inst_ack_1 : boolean;
  signal if_stmt_955_branch_ack_1 : boolean;
  signal type_cast_192_inst_req_1 : boolean;
  signal type_cast_634_inst_req_0 : boolean;
  signal type_cast_634_inst_ack_0 : boolean;
  signal type_cast_634_inst_req_1 : boolean;
  signal type_cast_153_inst_ack_0 : boolean;
  signal type_cast_634_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_648_inst_req_0 : boolean;
  signal type_cast_153_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_648_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_648_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_648_inst_ack_1 : boolean;
  signal if_stmt_955_branch_req_0 : boolean;
  signal type_cast_652_inst_req_0 : boolean;
  signal type_cast_652_inst_ack_0 : boolean;
  signal type_cast_652_inst_req_1 : boolean;
  signal type_cast_652_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_911_inst_ack_1 : boolean;
  signal ptr_deref_941_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_666_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_666_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_911_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_666_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_666_inst_ack_1 : boolean;
  signal ptr_deref_941_store_0_req_1 : boolean;
  signal type_cast_192_inst_ack_0 : boolean;
  signal type_cast_670_inst_req_0 : boolean;
  signal type_cast_670_inst_ack_0 : boolean;
  signal type_cast_670_inst_req_1 : boolean;
  signal type_cast_670_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_911_inst_ack_0 : boolean;
  signal ptr_deref_941_store_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_684_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_684_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_911_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_684_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_684_inst_ack_1 : boolean;
  signal ptr_deref_941_store_0_req_0 : boolean;
  signal type_cast_688_inst_req_0 : boolean;
  signal type_cast_688_inst_ack_0 : boolean;
  signal type_cast_192_inst_req_0 : boolean;
  signal type_cast_688_inst_req_1 : boolean;
  signal type_cast_688_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_702_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_702_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_702_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_702_inst_ack_1 : boolean;
  signal phi_stmt_189_ack_0 : boolean;
  signal type_cast_706_inst_req_0 : boolean;
  signal type_cast_706_inst_ack_0 : boolean;
  signal type_cast_706_inst_req_1 : boolean;
  signal type_cast_706_inst_ack_1 : boolean;
  signal type_cast_897_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_720_inst_req_0 : boolean;
  signal phi_stmt_80_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_720_inst_ack_0 : boolean;
  signal type_cast_897_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_720_inst_req_1 : boolean;
  signal phi_stmt_73_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_720_inst_ack_1 : boolean;
  signal type_cast_724_inst_req_0 : boolean;
  signal type_cast_724_inst_ack_0 : boolean;
  signal type_cast_724_inst_req_1 : boolean;
  signal type_cast_724_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_738_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_738_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_738_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_738_inst_ack_1 : boolean;
  signal type_cast_742_inst_req_0 : boolean;
  signal type_cast_742_inst_ack_0 : boolean;
  signal type_cast_742_inst_req_1 : boolean;
  signal type_cast_742_inst_ack_1 : boolean;
  signal ptr_deref_750_store_0_req_0 : boolean;
  signal ptr_deref_750_store_0_ack_0 : boolean;
  signal ptr_deref_750_store_0_req_1 : boolean;
  signal ptr_deref_750_store_0_ack_1 : boolean;
  signal if_stmt_764_branch_req_0 : boolean;
  signal if_stmt_764_branch_ack_1 : boolean;
  signal if_stmt_764_branch_ack_0 : boolean;
  signal array_obj_ref_804_index_offset_req_0 : boolean;
  signal array_obj_ref_804_index_offset_ack_0 : boolean;
  signal array_obj_ref_804_index_offset_req_1 : boolean;
  signal array_obj_ref_804_index_offset_ack_1 : boolean;
  signal addr_of_805_final_reg_req_0 : boolean;
  signal addr_of_805_final_reg_ack_0 : boolean;
  signal addr_of_805_final_reg_req_1 : boolean;
  signal addr_of_805_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_808_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_808_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_808_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_808_inst_ack_1 : boolean;
  signal type_cast_812_inst_req_0 : boolean;
  signal type_cast_812_inst_ack_0 : boolean;
  signal type_cast_812_inst_req_1 : boolean;
  signal type_cast_812_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_821_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_821_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_821_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_821_inst_ack_1 : boolean;
  signal type_cast_825_inst_req_0 : boolean;
  signal type_cast_825_inst_ack_0 : boolean;
  signal type_cast_825_inst_req_1 : boolean;
  signal type_cast_825_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_839_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_839_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_839_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_839_inst_ack_1 : boolean;
  signal type_cast_843_inst_req_0 : boolean;
  signal type_cast_843_inst_ack_0 : boolean;
  signal type_cast_843_inst_req_1 : boolean;
  signal type_cast_843_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_857_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_857_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_857_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_857_inst_ack_1 : boolean;
  signal type_cast_861_inst_req_0 : boolean;
  signal type_cast_861_inst_ack_0 : boolean;
  signal phi_stmt_270_req_0 : boolean;
  signal type_cast_280_inst_req_0 : boolean;
  signal type_cast_280_inst_ack_0 : boolean;
  signal type_cast_280_inst_req_1 : boolean;
  signal type_cast_280_inst_ack_1 : boolean;
  signal phi_stmt_277_req_0 : boolean;
  signal type_cast_276_inst_req_0 : boolean;
  signal type_cast_276_inst_ack_0 : boolean;
  signal type_cast_276_inst_req_1 : boolean;
  signal type_cast_276_inst_ack_1 : boolean;
  signal phi_stmt_270_req_1 : boolean;
  signal type_cast_282_inst_req_0 : boolean;
  signal type_cast_282_inst_ack_0 : boolean;
  signal type_cast_282_inst_req_1 : boolean;
  signal type_cast_282_inst_ack_1 : boolean;
  signal phi_stmt_277_req_1 : boolean;
  signal phi_stmt_270_ack_0 : boolean;
  signal phi_stmt_277_ack_0 : boolean;
  signal type_cast_322_inst_req_0 : boolean;
  signal type_cast_322_inst_ack_0 : boolean;
  signal type_cast_322_inst_req_1 : boolean;
  signal type_cast_322_inst_ack_1 : boolean;
  signal phi_stmt_319_req_0 : boolean;
  signal phi_stmt_319_ack_0 : boolean;
  signal phi_stmt_601_req_0 : boolean;
  signal type_cast_607_inst_req_0 : boolean;
  signal type_cast_607_inst_ack_0 : boolean;
  signal type_cast_607_inst_req_1 : boolean;
  signal type_cast_607_inst_ack_1 : boolean;
  signal phi_stmt_601_req_1 : boolean;
  signal phi_stmt_601_ack_0 : boolean;
  signal phi_stmt_792_req_0 : boolean;
  signal type_cast_798_inst_req_0 : boolean;
  signal type_cast_798_inst_ack_0 : boolean;
  signal type_cast_798_inst_req_1 : boolean;
  signal type_cast_798_inst_ack_1 : boolean;
  signal phi_stmt_792_req_1 : boolean;
  signal phi_stmt_792_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_0: Block -- control-path 
    signal testConfigure_CP_0_elements: BooleanArray(290 downto 0);
    -- 
  begin -- 
    testConfigure_CP_0_elements(0) <= testConfigure_CP_0_start;
    testConfigure_CP_0_symbol <= testConfigure_CP_0_elements(221);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (35) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/cr
      -- 
    rr_100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => ptr_deref_47_store_0_req_1); -- 
    cr_197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_62_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => testConfigure_CP_0_elements(1)); -- 
    cr_105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/rr
      -- 
    ca_106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => testConfigure_CP_0_elements(2)); -- 
    rr_114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_58_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/ra
      -- 
    ra_115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => testConfigure_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/ca
      -- 
    ca_120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => testConfigure_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/rr
      -- 
    rr_158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(5), ack => ptr_deref_47_store_0_req_0); -- 
    testConfigure_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(0) & testConfigure_CP_0_elements(4);
      gj_testConfigure_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/ra
      -- 
    ra_159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_47_store_0_ack_0, ack => testConfigure_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/ca
      -- 
    ca_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_47_store_0_ack_1, ack => testConfigure_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_update_start_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/cr
      -- 
    ra_179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_58_inst_ack_0, ack => testConfigure_CP_0_elements(8)); -- 
    cr_183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(8), ack => RPIPE_ConvTranspose_input_pipe_58_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/rr
      -- 
    ca_184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_58_inst_ack_1, ack => testConfigure_CP_0_elements(9)); -- 
    rr_192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(9), ack => type_cast_62_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/ra
      -- 
    ra_193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_62_inst_ack_0, ack => testConfigure_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/ca
      -- 
    ca_198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_62_inst_ack_1, ack => testConfigure_CP_0_elements(11)); -- 
    -- CP-element group 12:  branch  join  transition  place  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (10) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63__exit__
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64__entry__
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_32/R_cmp215_65_place
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_else_link/$entry
      -- 
    branch_req_206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(12), ack => if_stmt_64_branch_req_0); -- 
    testConfigure_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(7) & testConfigure_CP_0_elements(11);
      gj_testConfigure_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	242 
    -- CP-element group 13: 	243 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Update/cr
      -- CP-element group 13: 	 branch_block_stmt_32/if_stmt_64_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/if_stmt_64_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/$entry
      -- 
    if_choice_transition_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_64_branch_ack_1, ack => testConfigure_CP_0_elements(13)); -- 
    rr_2532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_160_inst_req_0); -- 
    cr_2537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_160_inst_req_1); -- 
    -- CP-element group 14:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	229 
    -- CP-element group 14: 	230 
    -- CP-element group 14: 	231 
    -- CP-element group 14:  members (22) 
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70__exit__
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/if_stmt_64_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/if_stmt_64_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/dummy
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/cr
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_64_branch_ack_0, ack => testConfigure_CP_0_elements(14)); -- 
    rr_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_85_inst_req_0); -- 
    cr_2470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_85_inst_req_1); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	237 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Sample/ra
      -- 
    ra_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => testConfigure_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	237 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	33 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Update/ca
      -- 
    ca_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => testConfigure_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	237 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	33 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_sample_complete
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Sample/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_0, ack => testConfigure_CP_0_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	237 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (11) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Update/ack
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_request/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_request/req
      -- 
    ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_1, ack => testConfigure_CP_0_elements(18)); -- 
    req_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(18), ack => addr_of_102_final_reg_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_request/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_request/ack
      -- 
    ack_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_0, ack => testConfigure_CP_0_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	237 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (28) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_complete/ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_root_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_address_resized
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_addr_resize/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_addr_resize/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_addr_resize/base_resize_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_addr_resize/base_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_plus_offset/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_plus_offset/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_plus_offset/sum_rename_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_base_plus_offset/sum_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_addrgen/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_addrgen/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_addrgen/root_register_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_word_addrgen/root_register_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/ptr_deref_105_Split/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/ptr_deref_105_Split/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/ptr_deref_105_Split/split_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/ptr_deref_105_Split/split_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/word_0/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/word_0/rr
      -- 
    ack_280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_1, ack => testConfigure_CP_0_elements(20)); -- 
    rr_318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(20), ack => ptr_deref_105_store_0_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	32 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Sample/word_access_start/word_0/ra
      -- 
    ra_319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_105_store_0_ack_0, ack => testConfigure_CP_0_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	237 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	33 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/word_0/ca
      -- 
    ca_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_105_store_0_ack_1, ack => testConfigure_CP_0_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	32 
    -- CP-element group 23: 	237 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/word_0/rr
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_sample_start_
      -- 
    rr_363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(23), ack => ptr_deref_122_load_0_req_0); -- 
    testConfigure_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(32) & testConfigure_CP_0_elements(237);
      gj_testConfigure_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Sample/word_access_start/word_0/ra
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_sample_completed_
      -- 
    ra_364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_122_load_0_ack_0, ack => testConfigure_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	237 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (12) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/ptr_deref_122_Merge/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/ptr_deref_122_Merge/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/ptr_deref_122_Merge/merge_req
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/ptr_deref_122_Merge/merge_ack
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Sample/rr
      -- 
    ca_375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_122_load_0_ack_1, ack => testConfigure_CP_0_elements(25)); -- 
    rr_388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(25), ack => type_cast_126_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Sample/ra
      -- 
    ra_389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => testConfigure_CP_0_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	237 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Update/ca
      -- 
    ca_394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => testConfigure_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	237 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_update_start_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Update/cr
      -- 
    ra_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_137_inst_ack_0, ack => testConfigure_CP_0_elements(28)); -- 
    cr_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(28), ack => RPIPE_ConvTranspose_input_pipe_137_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Sample/rr
      -- 
    ca_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_137_inst_ack_1, ack => testConfigure_CP_0_elements(29)); -- 
    rr_416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(29), ack => type_cast_141_inst_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Sample/ra
      -- 
    ra_417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_141_inst_ack_0, ack => testConfigure_CP_0_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	237 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Update/ca
      -- 
    ca_422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_141_inst_ack_1, ack => testConfigure_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  delay-element  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	21 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	23 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_ptr_deref_122_delay
      -- 
    -- Element group testConfigure_CP_0_elements(32) is a control-delay.
    cp_element_32_delay: control_delay_element  generic map(name => " 32_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(21), ack => testConfigure_CP_0_elements(32), clk => clk, reset =>reset);
    -- CP-element group 33:  branch  join  transition  place  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	17 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	27 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (10) 
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142__exit__
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143__entry__
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_dead_link/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_eval_test/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_eval_test/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_eval_test/branch_req
      -- CP-element group 33: 	 branch_block_stmt_32/R_cmp_144_place
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_if_link/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_143_else_link/$entry
      -- 
    branch_req_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => if_stmt_143_branch_req_0); -- 
    testConfigure_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(16) & testConfigure_CP_0_elements(17) & testConfigure_CP_0_elements(22) & testConfigure_CP_0_elements(27) & testConfigure_CP_0_elements(31);
      gj_testConfigure_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  place  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	222 
    -- CP-element group 34: 	223 
    -- CP-element group 34: 	225 
    -- CP-element group 34: 	226 
    -- CP-element group 34:  members (20) 
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/cr
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/if_stmt_143_if_link/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/if_stmt_143_if_link/if_choice_transition
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/cr
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/$entry
      -- 
    if_choice_transition_436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_143_branch_ack_1, ack => testConfigure_CP_0_elements(34)); -- 
    rr_2408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => type_cast_76_inst_req_0); -- 
    cr_2413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => type_cast_76_inst_req_1); -- 
    cr_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => type_cast_83_inst_req_1); -- 
    rr_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => type_cast_83_inst_req_0); -- 
    -- CP-element group 35:  fork  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	238 
    -- CP-element group 35: 	239 
    -- CP-element group 35:  members (12) 
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_143_else_link/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_143_else_link/else_choice_transition
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/cr
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- 
    else_choice_transition_440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_143_branch_ack_0, ack => testConfigure_CP_0_elements(35)); -- 
    cr_2506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => type_cast_153_inst_req_1); -- 
    rr_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => type_cast_153_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	249 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/word_0/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/word_0/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_171_store_0_ack_0, ack => testConfigure_CP_0_elements(36)); -- 
    -- CP-element group 37:  branch  transition  place  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	249 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (15) 
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179__exit__
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180__entry__
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/word_0/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/word_0/ca
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_dead_link/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_eval_test/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_eval_test/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_eval_test/branch_req
      -- CP-element group 37: 	 branch_block_stmt_32/R_cmp14210_181_place
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_if_link/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_180_else_link/$entry
      -- 
    ca_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_171_store_0_ack_1, ack => testConfigure_CP_0_elements(37)); -- 
    branch_req_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(37), ack => if_stmt_180_branch_req_0); -- 
    -- CP-element group 38:  transition  place  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	256 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_32/forx_xend_bbx_xnph207_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/if_stmt_180_if_link/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/if_stmt_180_if_link/if_choice_transition
      -- CP-element group 38: 	 branch_block_stmt_32/forx_xend_bbx_xnph207
      -- CP-element group 38: 	 branch_block_stmt_32/forx_xend_bbx_xnph207_PhiReq/$exit
      -- 
    if_choice_transition_508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_180_branch_ack_1, ack => testConfigure_CP_0_elements(38)); -- 
    -- CP-element group 39:  merge  transition  place  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	253 
    -- CP-element group 39:  members (14) 
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186__exit__
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16
      -- CP-element group 39: 	 branch_block_stmt_32/if_stmt_180_else_link/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/if_stmt_180_else_link/else_choice_transition
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xend_forx_xbody16x_xpreheader
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xend_forx_xbody16x_xpreheader_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xend_forx_xbody16x_xpreheader_PhiReq/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186_PhiAck/dummy
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186_PhiAck/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186_PhiAck/$entry
      -- CP-element group 39: 	 branch_block_stmt_32/merge_stmt_186_PhiReqMerge
      -- 
    else_choice_transition_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_180_branch_ack_0, ack => testConfigure_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	255 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Sample/ra
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_0, ack => testConfigure_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	255 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	59 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Update/ca
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_205_inst_ack_1, ack => testConfigure_CP_0_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	255 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	59 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_sample_complete
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Sample/ack
      -- 
    ack_557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_211_index_offset_ack_0, ack => testConfigure_CP_0_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	255 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (11) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_offset_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Update/ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_request/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_request/req
      -- 
    ack_562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_211_index_offset_ack_1, ack => testConfigure_CP_0_elements(43)); -- 
    req_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(43), ack => addr_of_212_final_reg_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_request/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_request/ack
      -- 
    ack_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_212_final_reg_ack_0, ack => testConfigure_CP_0_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	255 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	50 
    -- CP-element group 45:  members (19) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_complete/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_complete/ack
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_root_address_calculated
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_address_resized
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_addr_resize/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_addr_resize/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_addr_resize/base_resize_req
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_addr_resize/base_resize_ack
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_plus_offset/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_plus_offset/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_plus_offset/sum_rename_req
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_base_plus_offset/sum_rename_ack
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_addrgen/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_addrgen/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_addrgen/root_register_req
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_word_addrgen/root_register_ack
      -- 
    ack_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_212_final_reg_ack_1, ack => testConfigure_CP_0_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	255 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_update_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Update/cr
      -- 
    ra_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_215_inst_ack_0, ack => testConfigure_CP_0_elements(46)); -- 
    cr_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(46), ack => RPIPE_ConvTranspose_input_pipe_215_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Sample/rr
      -- 
    ca_591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_215_inst_ack_1, ack => testConfigure_CP_0_elements(47)); -- 
    rr_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(47), ack => type_cast_219_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Sample/ra
      -- 
    ra_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_0, ack => testConfigure_CP_0_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	255 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Update/ca
      -- 
    ca_605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_219_inst_ack_1, ack => testConfigure_CP_0_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/ptr_deref_222_Split/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/ptr_deref_222_Split/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/ptr_deref_222_Split/split_req
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/ptr_deref_222_Split/split_ack
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/word_0/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/word_0/rr
      -- 
    rr_643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(50), ack => ptr_deref_222_store_0_req_0); -- 
    testConfigure_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(45) & testConfigure_CP_0_elements(49);
      gj_testConfigure_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	58 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Sample/word_access_start/word_0/ra
      -- 
    ra_644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_store_0_ack_0, ack => testConfigure_CP_0_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	255 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	59 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/word_0/ca
      -- 
    ca_655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_store_0_ack_1, ack => testConfigure_CP_0_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	58 
    -- CP-element group 53: 	255 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/word_0/rr
      -- 
    rr_688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(53), ack => ptr_deref_239_load_0_req_0); -- 
    testConfigure_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(58) & testConfigure_CP_0_elements(255);
      gj_testConfigure_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Sample/word_access_start/word_0/ra
      -- 
    ra_689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_load_0_ack_0, ack => testConfigure_CP_0_elements(54)); -- 
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	255 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (12) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/ptr_deref_239_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/ptr_deref_239_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/ptr_deref_239_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/ptr_deref_239_Merge/merge_ack
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Sample/rr
      -- 
    ca_700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_load_0_ack_1, ack => testConfigure_CP_0_elements(55)); -- 
    rr_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => type_cast_243_inst_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Sample/ra
      -- 
    ra_714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_243_inst_ack_0, ack => testConfigure_CP_0_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	255 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Update/ca
      -- 
    ca_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_243_inst_ack_1, ack => testConfigure_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  delay-element  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	51 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	53 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_ptr_deref_239_delay
      -- 
    -- Element group testConfigure_CP_0_elements(58) is a control-delay.
    cp_element_58_delay: control_delay_element  generic map(name => " 58_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(51), ack => testConfigure_CP_0_elements(58), clk => clk, reset =>reset);
    -- CP-element group 59:  branch  join  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	41 
    -- CP-element group 59: 	42 
    -- CP-element group 59: 	52 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (10) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251__exit__
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252__entry__
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_32/R_cmp14_253_place
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/if_stmt_252_else_link/$entry
      -- 
    branch_req_728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(59), ack => if_stmt_252_branch_req_0); -- 
    testConfigure_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(41) & testConfigure_CP_0_elements(42) & testConfigure_CP_0_elements(52) & testConfigure_CP_0_elements(57);
      gj_testConfigure_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	250 
    -- CP-element group 60: 	251 
    -- CP-element group 60:  members (12) 
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/if_stmt_252_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_32/if_stmt_252_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Update/cr
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Sample/$entry
      -- 
    if_choice_transition_733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_252_branch_ack_1, ack => testConfigure_CP_0_elements(60)); -- 
    cr_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(60), ack => type_cast_192_inst_req_1); -- 
    rr_2601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(60), ack => type_cast_192_inst_req_0); -- 
    -- CP-element group 61:  merge  transition  place  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	256 
    -- CP-element group 61:  members (13) 
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258__exit__
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph207x_xloopexit_bbx_xnph207
      -- CP-element group 61: 	 branch_block_stmt_32/if_stmt_252_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/if_stmt_252_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_32/forx_xbody16_bbx_xnph207x_xloopexit
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph207x_xloopexit_bbx_xnph207_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258_PhiAck/dummy
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/merge_stmt_258_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_32/forx_xbody16_bbx_xnph207x_xloopexit_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/forx_xbody16_bbx_xnph207x_xloopexit_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph207x_xloopexit_bbx_xnph207_PhiReq/$exit
      -- 
    else_choice_transition_737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_252_branch_ack_0, ack => testConfigure_CP_0_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	256 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_update_start_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Sample/ra
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Update/cr
      -- 
    ra_751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_262_inst_ack_0, ack => testConfigure_CP_0_elements(62)); -- 
    cr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(62), ack => RPIPE_ConvTranspose_input_pipe_262_inst_req_1); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Update/ca
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Sample/rr
      -- 
    ca_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_262_inst_ack_1, ack => testConfigure_CP_0_elements(63)); -- 
    rr_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(63), ack => type_cast_266_inst_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Sample/ra
      -- 
    ra_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_0, ack => testConfigure_CP_0_elements(64)); -- 
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	256 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	257 
    -- CP-element group 65: 	258 
    -- CP-element group 65: 	259 
    -- CP-element group 65:  members (17) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267__exit__
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Update/ca
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_270/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Update/cr
      -- 
    ca_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_266_inst_ack_1, ack => testConfigure_CP_0_elements(65)); -- 
    rr_2674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(65), ack => type_cast_280_inst_req_0); -- 
    cr_2679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(65), ack => type_cast_280_inst_req_1); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	272 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_request/$exit
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_request/ack
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_sample_completed_
      -- 
    ack_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_287_final_reg_ack_0, ack => testConfigure_CP_0_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	272 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (28) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_complete/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_complete/ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_address_calculated
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_address_calculated
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_root_address_calculated
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_address_resized
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_addr_resize/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_addr_resize/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_addr_resize/base_resize_req
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_addr_resize/base_resize_ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_plus_offset/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_plus_offset/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_plus_offset/sum_rename_req
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_base_plus_offset/sum_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_addrgen/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_addrgen/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_addrgen/root_register_req
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_word_addrgen/root_register_ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/ptr_deref_290_Split/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/ptr_deref_290_Split/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/ptr_deref_290_Split/split_req
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/ptr_deref_290_Split/split_ack
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/word_0/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/word_0/rr
      -- 
    ack_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_287_final_reg_ack_1, ack => testConfigure_CP_0_elements(67)); -- 
    rr_850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(67), ack => ptr_deref_290_store_0_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/word_0/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Sample/word_access_start/word_0/ra
      -- 
    ra_851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_290_store_0_ack_0, ack => testConfigure_CP_0_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	272 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/word_0/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/word_0/ca
      -- 
    ca_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_290_store_0_ack_1, ack => testConfigure_CP_0_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	272 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_update_start_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Update/cr
      -- 
    ra_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_294_inst_ack_0, ack => testConfigure_CP_0_elements(70)); -- 
    cr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(70), ack => RPIPE_ConvTranspose_input_pipe_294_inst_req_1); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Sample/rr
      -- 
    ca_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_294_inst_ack_1, ack => testConfigure_CP_0_elements(71)); -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_298_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Sample/ra
      -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_298_inst_ack_0, ack => testConfigure_CP_0_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	272 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Update/ca
      -- 
    ca_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_298_inst_ack_1, ack => testConfigure_CP_0_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311__exit__
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312__entry__
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_32/R_exitcond9_313_place
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/if_stmt_312_else_link/$entry
      -- 
    branch_req_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(74), ack => if_stmt_312_branch_req_0); -- 
    testConfigure_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(69) & testConfigure_CP_0_elements(73);
      gj_testConfigure_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	273 
    -- CP-element group 75: 	274 
    -- CP-element group 75:  members (12) 
      -- CP-element group 75: 	 branch_block_stmt_32/if_stmt_312_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/if_stmt_312_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Update/cr
      -- 
    if_choice_transition_903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_312_branch_ack_1, ack => testConfigure_CP_0_elements(75)); -- 
    rr_2759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(75), ack => type_cast_322_inst_req_0); -- 
    cr_2764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(75), ack => type_cast_322_inst_req_1); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	262 
    -- CP-element group 76: 	263 
    -- CP-element group 76: 	265 
    -- CP-element group 76: 	266 
    -- CP-element group 76:  members (20) 
      -- CP-element group 76: 	 branch_block_stmt_32/if_stmt_312_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/if_stmt_312_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Update/cr
      -- 
    else_choice_transition_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_312_branch_ack_0, ack => testConfigure_CP_0_elements(76)); -- 
    rr_2700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => type_cast_276_inst_req_0); -- 
    cr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => type_cast_276_inst_req_1); -- 
    rr_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => type_cast_282_inst_req_0); -- 
    cr_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => type_cast_282_inst_req_1); -- 
    -- CP-element group 77:  join  fork  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	276 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	80 
    -- CP-element group 77: 	83 
    -- CP-element group 77: 	84 
    -- CP-element group 77: 	86 
    -- CP-element group 77: 	90 
    -- CP-element group 77: 	91 
    -- CP-element group 77: 	93 
    -- CP-element group 77: 	97 
    -- CP-element group 77: 	98 
    -- CP-element group 77: 	100 
    -- CP-element group 77: 	101 
    -- CP-element group 77: 	102 
    -- CP-element group 77: 	104 
    -- CP-element group 77: 	105 
    -- CP-element group 77: 	106 
    -- CP-element group 77: 	108 
    -- CP-element group 77: 	109 
    -- CP-element group 77: 	110 
    -- CP-element group 77: 	112 
    -- CP-element group 77: 	113 
    -- CP-element group 77: 	114 
    -- CP-element group 77: 	116 
    -- CP-element group 77: 	117 
    -- CP-element group 77: 	118 
    -- CP-element group 77: 	120 
    -- CP-element group 77: 	121 
    -- CP-element group 77: 	122 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	125 
    -- CP-element group 77: 	126 
    -- CP-element group 77: 	128 
    -- CP-element group 77:  members (295) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/STORE_padding_324_Split/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/STORE_padding_324_Split/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/STORE_padding_324_Split/split_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/STORE_padding_324_Split/split_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_word_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_address_resized
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_addr_resize/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_addr_resize/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_addr_resize/base_resize_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_addr_resize/base_resize_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_word_addrgen/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_word_addrgen/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_word_addrgen/root_register_req
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_word_addrgen/root_register_ack
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Sample/word_access_start/word_0/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/word_access_complete/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/word_access_complete/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/word_access_complete/word_0/cr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_Update/cr
      -- 
    cr_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => STORE_padding_324_store_0_req_1); -- 
    rr_933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => STORE_padding_324_store_0_req_0); -- 
    rr_953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => RPIPE_ConvTranspose_input_pipe_328_inst_req_0); -- 
    cr_972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_332_inst_req_1); -- 
    cr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_343_store_0_req_1); -- 
    cr_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_351_inst_req_1); -- 
    cr_1100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_362_store_0_req_1); -- 
    cr_1128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_370_inst_req_1); -- 
    cr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_381_store_0_req_1); -- 
    cr_1223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_394_load_0_req_1); -- 
    rr_1212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_394_load_0_req_0); -- 
    cr_1242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_398_inst_req_1); -- 
    cr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_410_load_0_req_1); -- 
    rr_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_410_load_0_req_0); -- 
    cr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_414_inst_req_1); -- 
    cr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_426_load_0_req_1); -- 
    rr_1340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_426_load_0_req_0); -- 
    cr_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_430_inst_req_1); -- 
    cr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_468_load_0_req_1); -- 
    rr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_468_load_0_req_0); -- 
    cr_1434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_472_inst_req_1); -- 
    cr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_484_load_0_req_1); -- 
    rr_1468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_484_load_0_req_0); -- 
    cr_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_488_inst_req_1); -- 
    cr_1543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_500_load_0_req_1); -- 
    rr_1532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_500_load_0_req_0); -- 
    cr_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_504_inst_req_1); -- 
    cr_1607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_516_load_0_req_1); -- 
    rr_1596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_516_load_0_req_0); -- 
    cr_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_520_inst_req_1); -- 
    testConfigure_CP_0_elements(77) <= testConfigure_CP_0_elements(276);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/word_access_start/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/word_access_start/word_0/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Sample/word_access_start/word_0/ra
      -- 
    ra_934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_324_store_0_ack_0, ack => testConfigure_CP_0_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	131 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Update/word_access_complete/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Update/word_access_complete/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/STORE_padding_324_Update/word_access_complete/word_0/ca
      -- 
    ca_945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_324_store_0_ack_1, ack => testConfigure_CP_0_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	77 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_update_start_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_Update/cr
      -- 
    ra_954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_328_inst_ack_0, ack => testConfigure_CP_0_elements(80)); -- 
    cr_958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(80), ack => RPIPE_ConvTranspose_input_pipe_328_inst_req_1); -- 
    -- CP-element group 81:  fork  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: 	87 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_328_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_Sample/rr
      -- 
    ca_959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_328_inst_ack_1, ack => testConfigure_CP_0_elements(81)); -- 
    rr_967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(81), ack => type_cast_332_inst_req_0); -- 
    rr_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(81), ack => RPIPE_ConvTranspose_input_pipe_347_inst_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_Sample/ra
      -- 
    ra_968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_332_inst_ack_0, ack => testConfigure_CP_0_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_332_Update/ca
      -- 
    ca_973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_332_inst_ack_1, ack => testConfigure_CP_0_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	77 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/ptr_deref_343_Split/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/ptr_deref_343_Split/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/ptr_deref_343_Split/split_req
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/ptr_deref_343_Split/split_ack
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/word_access_start/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/word_access_start/word_0/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/word_access_start/word_0/rr
      -- 
    rr_1011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => ptr_deref_343_store_0_req_0); -- 
    testConfigure_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(77) & testConfigure_CP_0_elements(83);
      gj_testConfigure_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	129 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/word_access_start/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/word_access_start/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Sample/word_access_start/word_0/ra
      -- 
    ra_1012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_343_store_0_ack_0, ack => testConfigure_CP_0_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	77 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	131 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Update/word_access_complete/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Update/word_access_complete/word_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_Update/word_access_complete/word_0/ca
      -- 
    ca_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_343_store_0_ack_1, ack => testConfigure_CP_0_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	81 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_update_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_Update/cr
      -- 
    ra_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_347_inst_ack_0, ack => testConfigure_CP_0_elements(87)); -- 
    cr_1036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(87), ack => RPIPE_ConvTranspose_input_pipe_347_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	94 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_347_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_Sample/rr
      -- 
    ca_1037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_347_inst_ack_1, ack => testConfigure_CP_0_elements(88)); -- 
    rr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(88), ack => type_cast_351_inst_req_0); -- 
    rr_1109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(88), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_Sample/ra
      -- 
    ra_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_351_inst_ack_0, ack => testConfigure_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	77 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_351_Update/ca
      -- 
    ca_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_351_inst_ack_1, ack => testConfigure_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	77 
    -- CP-element group 91: 	90 
    -- CP-element group 91: 	129 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/ptr_deref_362_Split/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/ptr_deref_362_Split/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/ptr_deref_362_Split/split_req
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/ptr_deref_362_Split/split_ack
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/word_access_start/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/word_access_start/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/word_access_start/word_0/rr
      -- 
    rr_1089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(91), ack => ptr_deref_362_store_0_req_0); -- 
    testConfigure_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(77) & testConfigure_CP_0_elements(90) & testConfigure_CP_0_elements(129);
      gj_testConfigure_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	130 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/word_access_start/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/word_access_start/word_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Sample/word_access_start/word_0/ra
      -- 
    ra_1090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_362_store_0_ack_0, ack => testConfigure_CP_0_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	77 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	131 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Update/word_access_complete/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Update/word_access_complete/word_0/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_Update/word_access_complete/word_0/ca
      -- 
    ca_1101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_362_store_0_ack_1, ack => testConfigure_CP_0_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	88 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_update_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_Update/cr
      -- 
    ra_1110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_0, ack => testConfigure_CP_0_elements(94)); -- 
    cr_1114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_1); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/RPIPE_ConvTranspose_input_pipe_366_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_sample_start_
      -- 
    ca_1115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_1, ack => testConfigure_CP_0_elements(95)); -- 
    rr_1123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(95), ack => type_cast_370_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_Sample/$exit
      -- 
    ra_1124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_0, ack => testConfigure_CP_0_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	77 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_370_update_completed_
      -- 
    ca_1129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_1, ack => testConfigure_CP_0_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	77 
    -- CP-element group 98: 	97 
    -- CP-element group 98: 	130 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/word_access_start/word_0/rr
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/word_access_start/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/word_access_start/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/ptr_deref_381_Split/split_ack
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/ptr_deref_381_Split/split_req
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/ptr_deref_381_Split/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/ptr_deref_381_Split/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/$entry
      -- 
    rr_1167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(98), ack => ptr_deref_381_store_0_req_0); -- 
    testConfigure_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(77) & testConfigure_CP_0_elements(97) & testConfigure_CP_0_elements(130);
      gj_testConfigure_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/word_access_start/word_0/ra
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/word_access_start/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Sample/$exit
      -- 
    ra_1168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_381_store_0_ack_0, ack => testConfigure_CP_0_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	77 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	131 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Update/word_access_complete/word_0/ca
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_381_Update/$exit
      -- 
    ca_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_381_store_0_ack_1, ack => testConfigure_CP_0_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	77 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Sample/word_access_start/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_sample_completed_
      -- 
    ra_1213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_394_load_0_ack_0, ack => testConfigure_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	77 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (12) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/ptr_deref_394_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/word_access_complete/word_0/ca
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/ptr_deref_394_Merge/merge_ack
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/ptr_deref_394_Merge/merge_req
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/ptr_deref_394_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/word_access_complete/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_394_update_completed_
      -- 
    ca_1224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_394_load_0_ack_1, ack => testConfigure_CP_0_elements(102)); -- 
    rr_1237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(102), ack => type_cast_398_inst_req_0); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_sample_completed_
      -- 
    ra_1238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_398_inst_ack_0, ack => testConfigure_CP_0_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	77 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	131 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_398_update_completed_
      -- 
    ca_1243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_398_inst_ack_1, ack => testConfigure_CP_0_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	77 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Sample/word_access_start/word_0/ra
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Sample/word_access_start/word_0/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Sample/word_access_start/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_sample_completed_
      -- 
    ra_1277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_410_load_0_ack_0, ack => testConfigure_CP_0_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	77 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (12) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/word_access_complete/word_0/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/ptr_deref_410_Merge/merge_ack
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/ptr_deref_410_Merge/merge_req
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/ptr_deref_410_Merge/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/ptr_deref_410_Merge/$entry
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/word_access_complete/word_0/ca
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/word_access_complete/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_Sample/rr
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_410_update_completed_
      -- 
    ca_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_410_load_0_ack_1, ack => testConfigure_CP_0_elements(106)); -- 
    rr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(106), ack => type_cast_414_inst_req_0); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_sample_completed_
      -- 
    ra_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_414_inst_ack_0, ack => testConfigure_CP_0_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	77 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	131 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_414_update_completed_
      -- 
    ca_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_414_inst_ack_1, ack => testConfigure_CP_0_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	77 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Sample/word_access_start/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Sample/word_access_start/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_sample_completed_
      -- 
    ra_1341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_426_load_0_ack_0, ack => testConfigure_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	77 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (12) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/word_access_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_Sample/rr
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/ptr_deref_426_Merge/merge_ack
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/ptr_deref_426_Merge/merge_req
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/ptr_deref_426_Merge/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/ptr_deref_426_Merge/$entry
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_426_update_completed_
      -- 
    ca_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_426_load_0_ack_1, ack => testConfigure_CP_0_elements(110)); -- 
    rr_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(110), ack => type_cast_430_inst_req_0); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_sample_completed_
      -- 
    ra_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_430_inst_ack_0, ack => testConfigure_CP_0_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	77 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	131 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_430_update_completed_
      -- 
    ca_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_430_inst_ack_1, ack => testConfigure_CP_0_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	77 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Sample/word_access_start/word_0/ra
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Sample/word_access_start/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Sample/word_access_start/$exit
      -- 
    ra_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_468_load_0_ack_0, ack => testConfigure_CP_0_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	77 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (12) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/ptr_deref_468_Merge/merge_ack
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/ptr_deref_468_Merge/merge_req
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/ptr_deref_468_Merge/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/ptr_deref_468_Merge/$entry
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/word_access_complete/word_0/ca
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/word_access_complete/word_0/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/word_access_complete/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_468_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_Sample/$entry
      -- 
    ca_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_468_load_0_ack_1, ack => testConfigure_CP_0_elements(114)); -- 
    rr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(114), ack => type_cast_472_inst_req_0); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_Sample/$exit
      -- 
    ra_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_472_inst_ack_0, ack => testConfigure_CP_0_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	77 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	131 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_472_Update/$exit
      -- 
    ca_1435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_472_inst_ack_1, ack => testConfigure_CP_0_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	77 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Sample/word_access_start/word_0/ra
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_sample_completed_
      -- 
    ra_1469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_484_load_0_ack_0, ack => testConfigure_CP_0_elements(117)); -- 
    -- CP-element group 118:  transition  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	77 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (12) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_Sample/rr
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/ptr_deref_484_Merge/merge_ack
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/ptr_deref_484_Merge/merge_req
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/ptr_deref_484_Merge/$exit
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_484_Update/ptr_deref_484_Merge/$entry
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_Sample/$entry
      -- 
    ca_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_484_load_0_ack_1, ack => testConfigure_CP_0_elements(118)); -- 
    rr_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(118), ack => type_cast_488_inst_req_0); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_Sample/$exit
      -- 
    ra_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_488_inst_ack_0, ack => testConfigure_CP_0_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	77 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	131 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_488_update_completed_
      -- 
    ca_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_488_inst_ack_1, ack => testConfigure_CP_0_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	77 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Sample/word_access_start/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Sample/word_access_start/word_0/ra
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Sample/word_access_start/word_0/$exit
      -- 
    ra_1533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_500_load_0_ack_0, ack => testConfigure_CP_0_elements(121)); -- 
    -- CP-element group 122:  transition  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	77 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (12) 
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/ptr_deref_500_Merge/merge_req
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/ptr_deref_500_Merge/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/ptr_deref_500_Merge/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/word_access_complete/word_0/ca
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/word_access_complete/word_0/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/word_access_complete/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_500_Update/ptr_deref_500_Merge/merge_ack
      -- 
    ca_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_500_load_0_ack_1, ack => testConfigure_CP_0_elements(122)); -- 
    rr_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(122), ack => type_cast_504_inst_req_0); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_Sample/ra
      -- 
    ra_1558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_0, ack => testConfigure_CP_0_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	131 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_504_Update/ca
      -- 
    ca_1563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_1, ack => testConfigure_CP_0_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	77 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Sample/word_access_start/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Sample/word_access_start/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Sample/word_access_start/word_0/ra
      -- 
    ra_1597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_516_load_0_ack_0, ack => testConfigure_CP_0_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	77 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (12) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/word_access_complete/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/word_access_complete/word_0/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/word_access_complete/word_0/ca
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/ptr_deref_516_Merge/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/ptr_deref_516_Merge/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/ptr_deref_516_Merge/merge_req
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_516_Update/ptr_deref_516_Merge/merge_ack
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_Sample/rr
      -- 
    ca_1608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_516_load_0_ack_1, ack => testConfigure_CP_0_elements(126)); -- 
    rr_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(126), ack => type_cast_520_inst_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_Sample/ra
      -- 
    ra_1622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_0, ack => testConfigure_CP_0_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	77 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	131 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/type_cast_520_Update/ca
      -- 
    ca_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_520_inst_ack_1, ack => testConfigure_CP_0_elements(128)); -- 
    -- CP-element group 129:  transition  delay-element  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	85 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	91 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_343_ptr_deref_362_delay
      -- 
    -- Element group testConfigure_CP_0_elements(129) is a control-delay.
    cp_element_129_delay: control_delay_element  generic map(name => " 129_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(85), ack => testConfigure_CP_0_elements(129), clk => clk, reset =>reset);
    -- CP-element group 130:  transition  delay-element  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	92 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	98 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/ptr_deref_362_ptr_deref_381_delay
      -- 
    -- Element group testConfigure_CP_0_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(92), ack => testConfigure_CP_0_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  branch  join  transition  place  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	79 
    -- CP-element group 131: 	86 
    -- CP-element group 131: 	93 
    -- CP-element group 131: 	100 
    -- CP-element group 131: 	104 
    -- CP-element group 131: 	108 
    -- CP-element group 131: 	112 
    -- CP-element group 131: 	116 
    -- CP-element group 131: 	120 
    -- CP-element group 131: 	124 
    -- CP-element group 131: 	128 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (10) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557__exit__
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_558__entry__
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_558_dead_link/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_558_eval_test/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_558_eval_test/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_558_eval_test/branch_req
      -- CP-element group 131: 	 branch_block_stmt_32/R_cmp74199_559_place
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_558_if_link/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/if_stmt_558_else_link/$entry
      -- 
    branch_req_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => if_stmt_558_branch_req_0); -- 
    testConfigure_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(79) & testConfigure_CP_0_elements(86) & testConfigure_CP_0_elements(93) & testConfigure_CP_0_elements(100) & testConfigure_CP_0_elements(104) & testConfigure_CP_0_elements(108) & testConfigure_CP_0_elements(112) & testConfigure_CP_0_elements(116) & testConfigure_CP_0_elements(120) & testConfigure_CP_0_elements(124) & testConfigure_CP_0_elements(128);
      gj_testConfigure_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  merge  transition  place  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	278 
    -- CP-element group 132:  members (18) 
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_579__exit__
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_585_to_assign_stmt_598__entry__
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_585_to_assign_stmt_598__exit__
      -- CP-element group 132: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76
      -- CP-element group 132: 	 branch_block_stmt_32/if_stmt_558_if_link/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/if_stmt_558_if_link/if_choice_transition
      -- CP-element group 132: 	 branch_block_stmt_32/forx_xend39_bbx_xnph201
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_585_to_assign_stmt_598/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_585_to_assign_stmt_598/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/forx_xend39_bbx_xnph201_PhiReq/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/forx_xend39_bbx_xnph201_PhiReq/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_579_PhiReqMerge
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_579_PhiAck/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_579_PhiAck/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/merge_stmt_579_PhiAck/dummy
      -- CP-element group 132: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76_PhiReq/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76_PhiReq/phi_stmt_601/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/$entry
      -- 
    if_choice_transition_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_558_branch_ack_1, ack => testConfigure_CP_0_elements(132)); -- 
    -- CP-element group 133:  transition  place  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	277 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_32/if_stmt_558_else_link/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/if_stmt_558_else_link/else_choice_transition
      -- CP-element group 133: 	 branch_block_stmt_32/forx_xend39_forx_xcond128x_xpreheader
      -- CP-element group 133: 	 branch_block_stmt_32/forx_xend39_forx_xcond128x_xpreheader_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_32/forx_xend39_forx_xcond128x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_1646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_558_branch_ack_0, ack => testConfigure_CP_0_elements(133)); -- 
    -- CP-element group 134:  merge  transition  place  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	277 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	284 
    -- CP-element group 134:  members (18) 
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_770__exit__
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_776_to_assign_stmt_789__entry__
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_776_to_assign_stmt_789__exit__
      -- CP-element group 134: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135
      -- CP-element group 134: 	 branch_block_stmt_32/if_stmt_573_if_link/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/if_stmt_573_if_link/if_choice_transition
      -- CP-element group 134: 	 branch_block_stmt_32/forx_xcond128x_xpreheader_bbx_xnph
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_776_to_assign_stmt_789/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_776_to_assign_stmt_789/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/forx_xcond128x_xpreheader_bbx_xnph_PhiReq/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/forx_xcond128x_xpreheader_bbx_xnph_PhiReq/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_770_PhiReqMerge
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_770_PhiAck/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_770_PhiAck/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/merge_stmt_770_PhiAck/dummy
      -- CP-element group 134: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135_PhiReq/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135_PhiReq/phi_stmt_792/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/$entry
      -- 
    if_choice_transition_1664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_573_branch_ack_1, ack => testConfigure_CP_0_elements(134)); -- 
    -- CP-element group 135:  transition  place  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	277 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	290 
    -- CP-element group 135:  members (5) 
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_573_else_link/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/if_stmt_573_else_link/else_choice_transition
      -- CP-element group 135: 	 branch_block_stmt_32/forx_xcond128x_xpreheader_forx_xend189
      -- CP-element group 135: 	 branch_block_stmt_32/forx_xcond128x_xpreheader_forx_xend189_PhiReq/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/forx_xcond128x_xpreheader_forx_xend189_PhiReq/$exit
      -- 
    else_choice_transition_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_573_branch_ack_0, ack => testConfigure_CP_0_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	283 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	175 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_sample_complete
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_Sample/ack
      -- 
    ack_1702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_613_index_offset_ack_0, ack => testConfigure_CP_0_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	283 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (11) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_root_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_offset_calculated
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_Update/ack
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_base_plus_offset/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_base_plus_offset/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_base_plus_offset/sum_rename_req
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_base_plus_offset/sum_rename_ack
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_request/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_request/req
      -- 
    ack_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_613_index_offset_ack_1, ack => testConfigure_CP_0_elements(137)); -- 
    req_1716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(137), ack => addr_of_614_final_reg_req_0); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_request/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_request/ack
      -- 
    ack_1717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_614_final_reg_ack_0, ack => testConfigure_CP_0_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	283 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	172 
    -- CP-element group 139:  members (19) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_complete/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_complete/ack
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_word_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_address_resized
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_addr_resize/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_addr_resize/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_addr_resize/base_resize_req
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_addr_resize/base_resize_ack
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_plus_offset/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_plus_offset/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_plus_offset/sum_rename_req
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_base_plus_offset/sum_rename_ack
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_word_addrgen/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_word_addrgen/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_word_addrgen/root_register_req
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_word_addrgen/root_register_ack
      -- 
    ack_1722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_614_final_reg_ack_1, ack => testConfigure_CP_0_elements(139)); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	283 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (6) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_update_start_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_Sample/ra
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_Update/cr
      -- 
    ra_1731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_617_inst_ack_0, ack => testConfigure_CP_0_elements(140)); -- 
    cr_1735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(140), ack => RPIPE_ConvTranspose_input_pipe_617_inst_req_1); -- 
    -- CP-element group 141:  fork  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141: 	144 
    -- CP-element group 141:  members (9) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_Update/ca
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_Sample/rr
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_Sample/rr
      -- 
    ca_1736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_617_inst_ack_1, ack => testConfigure_CP_0_elements(141)); -- 
    rr_1744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(141), ack => type_cast_621_inst_req_0); -- 
    rr_1758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(141), ack => RPIPE_ConvTranspose_input_pipe_630_inst_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_Sample/ra
      -- 
    ra_1745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_621_inst_ack_0, ack => testConfigure_CP_0_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	283 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	172 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_Update/ca
      -- 
    ca_1750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_621_inst_ack_1, ack => testConfigure_CP_0_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	141 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (6) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_update_start_
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_Sample/ra
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_Update/cr
      -- 
    ra_1759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_630_inst_ack_0, ack => testConfigure_CP_0_elements(144)); -- 
    cr_1763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(144), ack => RPIPE_ConvTranspose_input_pipe_630_inst_req_1); -- 
    -- CP-element group 145:  fork  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145: 	148 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_630_Update/ca
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_Sample/rr
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_Sample/rr
      -- 
    ca_1764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_630_inst_ack_1, ack => testConfigure_CP_0_elements(145)); -- 
    rr_1772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(145), ack => type_cast_634_inst_req_0); -- 
    rr_1786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(145), ack => RPIPE_ConvTranspose_input_pipe_648_inst_req_0); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_Sample/ra
      -- 
    ra_1773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_634_inst_ack_0, ack => testConfigure_CP_0_elements(146)); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	283 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	172 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_Update/ca
      -- 
    ca_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_634_inst_ack_1, ack => testConfigure_CP_0_elements(147)); -- 
    -- CP-element group 148:  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	145 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (6) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_update_start_
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_Sample/ra
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_Update/cr
      -- 
    ra_1787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_648_inst_ack_0, ack => testConfigure_CP_0_elements(148)); -- 
    cr_1791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(148), ack => RPIPE_ConvTranspose_input_pipe_648_inst_req_1); -- 
    -- CP-element group 149:  fork  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149: 	152 
    -- CP-element group 149:  members (9) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_648_Update/ca
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_Sample/rr
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_Sample/rr
      -- 
    ca_1792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_648_inst_ack_1, ack => testConfigure_CP_0_elements(149)); -- 
    rr_1800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(149), ack => type_cast_652_inst_req_0); -- 
    rr_1814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(149), ack => RPIPE_ConvTranspose_input_pipe_666_inst_req_0); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_Sample/ra
      -- 
    ra_1801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_0, ack => testConfigure_CP_0_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	283 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	172 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_Update/ca
      -- 
    ca_1806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_652_inst_ack_1, ack => testConfigure_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	149 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_update_start_
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_Update/cr
      -- 
    ra_1815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_666_inst_ack_0, ack => testConfigure_CP_0_elements(152)); -- 
    cr_1819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(152), ack => RPIPE_ConvTranspose_input_pipe_666_inst_req_1); -- 
    -- CP-element group 153:  fork  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	156 
    -- CP-element group 153:  members (9) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_666_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_Sample/rr
      -- 
    ca_1820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_666_inst_ack_1, ack => testConfigure_CP_0_elements(153)); -- 
    rr_1828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(153), ack => type_cast_670_inst_req_0); -- 
    rr_1842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(153), ack => RPIPE_ConvTranspose_input_pipe_684_inst_req_0); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_Sample/ra
      -- 
    ra_1829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_670_inst_ack_0, ack => testConfigure_CP_0_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	283 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	172 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_Update/ca
      -- 
    ca_1834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_670_inst_ack_1, ack => testConfigure_CP_0_elements(155)); -- 
    -- CP-element group 156:  transition  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	153 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (6) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_update_start_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_Update/cr
      -- 
    ra_1843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_684_inst_ack_0, ack => testConfigure_CP_0_elements(156)); -- 
    cr_1847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(156), ack => RPIPE_ConvTranspose_input_pipe_684_inst_req_1); -- 
    -- CP-element group 157:  fork  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: 	160 
    -- CP-element group 157:  members (9) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_684_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_Sample/rr
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_Sample/rr
      -- 
    ca_1848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_684_inst_ack_1, ack => testConfigure_CP_0_elements(157)); -- 
    rr_1856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(157), ack => type_cast_688_inst_req_0); -- 
    rr_1870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(157), ack => RPIPE_ConvTranspose_input_pipe_702_inst_req_0); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_Sample/ra
      -- 
    ra_1857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_0, ack => testConfigure_CP_0_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	283 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	172 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_Update/ca
      -- 
    ca_1862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_688_inst_ack_1, ack => testConfigure_CP_0_elements(159)); -- 
    -- CP-element group 160:  transition  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	157 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (6) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_update_start_
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_Sample/ra
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_Update/cr
      -- 
    ra_1871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_702_inst_ack_0, ack => testConfigure_CP_0_elements(160)); -- 
    cr_1875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(160), ack => RPIPE_ConvTranspose_input_pipe_702_inst_req_1); -- 
    -- CP-element group 161:  fork  transition  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: 	164 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_702_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_Sample/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_Sample/rr
      -- 
    ca_1876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_702_inst_ack_1, ack => testConfigure_CP_0_elements(161)); -- 
    rr_1884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(161), ack => type_cast_706_inst_req_0); -- 
    rr_1898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(161), ack => RPIPE_ConvTranspose_input_pipe_720_inst_req_0); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_Sample/ra
      -- 
    ra_1885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_706_inst_ack_0, ack => testConfigure_CP_0_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	283 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	172 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_Update/ca
      -- 
    ca_1890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_706_inst_ack_1, ack => testConfigure_CP_0_elements(163)); -- 
    -- CP-element group 164:  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	161 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_update_start_
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_Sample/ra
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_Update/cr
      -- 
    ra_1899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_720_inst_ack_0, ack => testConfigure_CP_0_elements(164)); -- 
    cr_1903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(164), ack => RPIPE_ConvTranspose_input_pipe_720_inst_req_1); -- 
    -- CP-element group 165:  fork  transition  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	168 
    -- CP-element group 165:  members (9) 
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_720_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_Sample/rr
      -- 
    ca_1904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_720_inst_ack_1, ack => testConfigure_CP_0_elements(165)); -- 
    rr_1912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(165), ack => type_cast_724_inst_req_0); -- 
    rr_1926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(165), ack => RPIPE_ConvTranspose_input_pipe_738_inst_req_0); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_Sample/ra
      -- 
    ra_1913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_724_inst_ack_0, ack => testConfigure_CP_0_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	283 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	172 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_Update/ca
      -- 
    ca_1918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_724_inst_ack_1, ack => testConfigure_CP_0_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	165 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_update_start_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_Sample/ra
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_Update/cr
      -- 
    ra_1927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_738_inst_ack_0, ack => testConfigure_CP_0_elements(168)); -- 
    cr_1931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(168), ack => RPIPE_ConvTranspose_input_pipe_738_inst_req_1); -- 
    -- CP-element group 169:  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (6) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_738_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_Sample/rr
      -- 
    ca_1932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_738_inst_ack_1, ack => testConfigure_CP_0_elements(169)); -- 
    rr_1940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(169), ack => type_cast_742_inst_req_0); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_Sample/ra
      -- 
    ra_1941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_742_inst_ack_0, ack => testConfigure_CP_0_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	283 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_Update/ca
      -- 
    ca_1946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_742_inst_ack_1, ack => testConfigure_CP_0_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	139 
    -- CP-element group 172: 	143 
    -- CP-element group 172: 	147 
    -- CP-element group 172: 	151 
    -- CP-element group 172: 	155 
    -- CP-element group 172: 	159 
    -- CP-element group 172: 	163 
    -- CP-element group 172: 	167 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (9) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/ptr_deref_750_Split/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/ptr_deref_750_Split/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/ptr_deref_750_Split/split_req
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/ptr_deref_750_Split/split_ack
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/word_access_start/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/word_access_start/word_0/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/word_access_start/word_0/rr
      -- 
    rr_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(172), ack => ptr_deref_750_store_0_req_0); -- 
    testConfigure_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(139) & testConfigure_CP_0_elements(143) & testConfigure_CP_0_elements(147) & testConfigure_CP_0_elements(151) & testConfigure_CP_0_elements(155) & testConfigure_CP_0_elements(159) & testConfigure_CP_0_elements(163) & testConfigure_CP_0_elements(167) & testConfigure_CP_0_elements(171);
      gj_testConfigure_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (5) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/word_access_start/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/word_access_start/word_0/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Sample/word_access_start/word_0/ra
      -- 
    ra_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_750_store_0_ack_0, ack => testConfigure_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	283 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (5) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Update/word_access_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Update/word_access_complete/word_0/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Update/word_access_complete/word_0/ca
      -- 
    ca_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_750_store_0_ack_1, ack => testConfigure_CP_0_elements(174)); -- 
    -- CP-element group 175:  branch  join  transition  place  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	136 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (10) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763__exit__
      -- CP-element group 175: 	 branch_block_stmt_32/if_stmt_764__entry__
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/if_stmt_764_dead_link/$entry
      -- CP-element group 175: 	 branch_block_stmt_32/if_stmt_764_eval_test/$entry
      -- CP-element group 175: 	 branch_block_stmt_32/if_stmt_764_eval_test/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/if_stmt_764_eval_test/branch_req
      -- CP-element group 175: 	 branch_block_stmt_32/R_exitcond_765_place
      -- CP-element group 175: 	 branch_block_stmt_32/if_stmt_764_if_link/$entry
      -- CP-element group 175: 	 branch_block_stmt_32/if_stmt_764_else_link/$entry
      -- 
    branch_req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => if_stmt_764_branch_req_0); -- 
    testConfigure_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(136) & testConfigure_CP_0_elements(174);
      gj_testConfigure_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  merge  transition  place  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	277 
    -- CP-element group 176:  members (13) 
      -- CP-element group 176: 	 branch_block_stmt_32/merge_stmt_564__exit__
      -- CP-element group 176: 	 branch_block_stmt_32/forx_xcond128x_xpreheaderx_xloopexit_forx_xcond128x_xpreheader
      -- CP-element group 176: 	 branch_block_stmt_32/if_stmt_764_if_link/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/if_stmt_764_if_link/if_choice_transition
      -- CP-element group 176: 	 branch_block_stmt_32/forx_xbody76_forx_xcond128x_xpreheaderx_xloopexit
      -- CP-element group 176: 	 branch_block_stmt_32/forx_xbody76_forx_xcond128x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 176: 	 branch_block_stmt_32/forx_xbody76_forx_xcond128x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/merge_stmt_564_PhiReqMerge
      -- CP-element group 176: 	 branch_block_stmt_32/merge_stmt_564_PhiAck/$entry
      -- CP-element group 176: 	 branch_block_stmt_32/merge_stmt_564_PhiAck/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/merge_stmt_564_PhiAck/dummy
      -- CP-element group 176: 	 branch_block_stmt_32/forx_xcond128x_xpreheaderx_xloopexit_forx_xcond128x_xpreheader_PhiReq/$entry
      -- CP-element group 176: 	 branch_block_stmt_32/forx_xcond128x_xpreheaderx_xloopexit_forx_xcond128x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_2009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_764_branch_ack_1, ack => testConfigure_CP_0_elements(176)); -- 
    -- CP-element group 177:  fork  transition  place  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	279 
    -- CP-element group 177: 	280 
    -- CP-element group 177:  members (12) 
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_764_else_link/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/if_stmt_764_else_link/else_choice_transition
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/Sample/rr
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_764_branch_ack_0, ack => testConfigure_CP_0_elements(177)); -- 
    rr_2836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(177), ack => type_cast_607_inst_req_0); -- 
    cr_2841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(177), ack => type_cast_607_inst_req_1); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	289 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	217 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_sample_complete
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_Sample/ack
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_804_index_offset_ack_0, ack => testConfigure_CP_0_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	289 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (11) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_root_address_calculated
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_offset_calculated
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_Update/ack
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_base_plus_offset/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_base_plus_offset/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_base_plus_offset/sum_rename_req
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_base_plus_offset/sum_rename_ack
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_request/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_request/req
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_804_index_offset_ack_1, ack => testConfigure_CP_0_elements(179)); -- 
    req_2061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => addr_of_805_final_reg_req_0); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_request/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_request/ack
      -- 
    ack_2062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_805_final_reg_ack_0, ack => testConfigure_CP_0_elements(180)); -- 
    -- CP-element group 181:  fork  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	289 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	214 
    -- CP-element group 181:  members (19) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_address_calculated
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_word_address_calculated
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_root_address_calculated
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_address_resized
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_addr_resize/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_addr_resize/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_word_addrgen/root_register_ack
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_word_addrgen/root_register_req
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_word_addrgen/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_word_addrgen/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_plus_offset/sum_rename_ack
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_plus_offset/sum_rename_req
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_plus_offset/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_plus_offset/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_addr_resize/base_resize_ack
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_base_addr_resize/base_resize_req
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_complete/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_complete/ack
      -- 
    ack_2067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_805_final_reg_ack_1, ack => testConfigure_CP_0_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	289 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (6) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_update_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_Sample/ra
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_Update/cr
      -- 
    ra_2076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_808_inst_ack_0, ack => testConfigure_CP_0_elements(182)); -- 
    cr_2080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(182), ack => RPIPE_ConvTranspose_input_pipe_808_inst_req_1); -- 
    -- CP-element group 183:  fork  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183: 	186 
    -- CP-element group 183:  members (9) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_Update/ca
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_Sample/rr
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_Sample/rr
      -- 
    ca_2081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_808_inst_ack_1, ack => testConfigure_CP_0_elements(183)); -- 
    rr_2089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => type_cast_812_inst_req_0); -- 
    rr_2103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => RPIPE_ConvTranspose_input_pipe_821_inst_req_0); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_Sample/ra
      -- 
    ra_2090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_812_inst_ack_0, ack => testConfigure_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	289 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	214 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_Update/ca
      -- 
    ca_2095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_812_inst_ack_1, ack => testConfigure_CP_0_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	183 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_update_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_Update/cr
      -- 
    ra_2104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_821_inst_ack_0, ack => testConfigure_CP_0_elements(186)); -- 
    cr_2108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(186), ack => RPIPE_ConvTranspose_input_pipe_821_inst_req_1); -- 
    -- CP-element group 187:  fork  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	190 
    -- CP-element group 187:  members (9) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_821_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_Sample/rr
      -- 
    ca_2109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_821_inst_ack_1, ack => testConfigure_CP_0_elements(187)); -- 
    rr_2117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => type_cast_825_inst_req_0); -- 
    rr_2131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => RPIPE_ConvTranspose_input_pipe_839_inst_req_0); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_Sample/ra
      -- 
    ra_2118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_825_inst_ack_0, ack => testConfigure_CP_0_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	289 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	214 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_Update/ca
      -- 
    ca_2123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_825_inst_ack_1, ack => testConfigure_CP_0_elements(189)); -- 
    -- CP-element group 190:  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	187 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (6) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_update_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_Sample/ra
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_Update/cr
      -- 
    ra_2132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_839_inst_ack_0, ack => testConfigure_CP_0_elements(190)); -- 
    cr_2136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(190), ack => RPIPE_ConvTranspose_input_pipe_839_inst_req_1); -- 
    -- CP-element group 191:  fork  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191: 	194 
    -- CP-element group 191:  members (9) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_839_Update/ca
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_Sample/rr
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_Sample/rr
      -- 
    ca_2137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_839_inst_ack_1, ack => testConfigure_CP_0_elements(191)); -- 
    rr_2145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => type_cast_843_inst_req_0); -- 
    rr_2159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => RPIPE_ConvTranspose_input_pipe_857_inst_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_Sample/ra
      -- 
    ra_2146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_0, ack => testConfigure_CP_0_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	289 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	214 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_Update/ca
      -- 
    ca_2151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_843_inst_ack_1, ack => testConfigure_CP_0_elements(193)); -- 
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	191 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_update_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_Update/cr
      -- 
    ra_2160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_857_inst_ack_0, ack => testConfigure_CP_0_elements(194)); -- 
    cr_2164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(194), ack => RPIPE_ConvTranspose_input_pipe_857_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195: 	198 
    -- CP-element group 195:  members (9) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_857_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_Sample/rr
      -- 
    ca_2165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_857_inst_ack_1, ack => testConfigure_CP_0_elements(195)); -- 
    rr_2173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => type_cast_861_inst_req_0); -- 
    rr_2187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => RPIPE_ConvTranspose_input_pipe_875_inst_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_Sample/ra
      -- 
    ra_2174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_0, ack => testConfigure_CP_0_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	289 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	214 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_Update/ca
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_update_completed_
      -- 
    ca_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_861_inst_ack_1, ack => testConfigure_CP_0_elements(197)); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	195 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_update_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_Update/cr
      -- 
    ra_2188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_875_inst_ack_0, ack => testConfigure_CP_0_elements(198)); -- 
    cr_2192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(198), ack => RPIPE_ConvTranspose_input_pipe_875_inst_req_1); -- 
    -- CP-element group 199:  fork  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: 	202 
    -- CP-element group 199:  members (9) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_875_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_sample_start_
      -- 
    ca_2193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_875_inst_ack_1, ack => testConfigure_CP_0_elements(199)); -- 
    rr_2201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => type_cast_879_inst_req_0); -- 
    rr_2215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => RPIPE_ConvTranspose_input_pipe_893_inst_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_Sample/ra
      -- 
    ra_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_879_inst_ack_0, ack => testConfigure_CP_0_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	289 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	214 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_Update/ca
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_Update/$exit
      -- 
    ca_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_879_inst_ack_1, ack => testConfigure_CP_0_elements(201)); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	199 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_Update/cr
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_update_start_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_sample_completed_
      -- 
    ra_2216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_893_inst_ack_0, ack => testConfigure_CP_0_elements(202)); -- 
    cr_2220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(202), ack => RPIPE_ConvTranspose_input_pipe_893_inst_req_1); -- 
    -- CP-element group 203:  fork  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203: 	206 
    -- CP-element group 203:  members (9) 
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_Update/ca
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_Sample/rr
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_893_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_Sample/rr
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_sample_start_
      -- 
    ca_2221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_893_inst_ack_1, ack => testConfigure_CP_0_elements(203)); -- 
    rr_2229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => type_cast_897_inst_req_0); -- 
    rr_2243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => RPIPE_ConvTranspose_input_pipe_911_inst_req_0); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_Sample/ra
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_Sample/$exit
      -- 
    ra_2230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_0, ack => testConfigure_CP_0_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	289 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	214 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_Update/ca
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_Update/$exit
      -- 
    ca_2235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_1, ack => testConfigure_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	203 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (6) 
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_Update/cr
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_Sample/ra
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_update_start_
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_sample_completed_
      -- 
    ra_2244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_911_inst_ack_0, ack => testConfigure_CP_0_elements(206)); -- 
    cr_2248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(206), ack => RPIPE_ConvTranspose_input_pipe_911_inst_req_1); -- 
    -- CP-element group 207:  fork  transition  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207: 	210 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_Update/ca
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_911_update_completed_
      -- 
    ca_2249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_911_inst_ack_1, ack => testConfigure_CP_0_elements(207)); -- 
    rr_2257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(207), ack => type_cast_915_inst_req_0); -- 
    rr_2271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(207), ack => RPIPE_ConvTranspose_input_pipe_929_inst_req_0); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_Sample/ra
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_sample_completed_
      -- 
    ra_2258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_0, ack => testConfigure_CP_0_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	289 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	214 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_Update/ca
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_update_completed_
      -- 
    ca_2263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_1, ack => testConfigure_CP_0_elements(209)); -- 
    -- CP-element group 210:  transition  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	207 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (6) 
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_Sample/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_Sample/ra
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_Update/cr
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_sample_completed_
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_update_start_
      -- 
    ra_2272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_929_inst_ack_0, ack => testConfigure_CP_0_elements(210)); -- 
    cr_2276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(210), ack => RPIPE_ConvTranspose_input_pipe_929_inst_req_1); -- 
    -- CP-element group 211:  transition  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211:  members (6) 
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_update_completed_
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_Update/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_929_Update/ca
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_Sample/rr
      -- 
    ca_2277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_929_inst_ack_1, ack => testConfigure_CP_0_elements(211)); -- 
    rr_2285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_933_inst_req_0); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_Sample/ra
      -- 
    ra_2286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_933_inst_ack_0, ack => testConfigure_CP_0_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	289 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_Update/ca
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_Update/$exit
      -- 
    ca_2291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_933_inst_ack_1, ack => testConfigure_CP_0_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	181 
    -- CP-element group 214: 	185 
    -- CP-element group 214: 	189 
    -- CP-element group 214: 	193 
    -- CP-element group 214: 	197 
    -- CP-element group 214: 	201 
    -- CP-element group 214: 	205 
    -- CP-element group 214: 	209 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (9) 
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/word_access_start/word_0/rr
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/word_access_start/word_0/$entry
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/word_access_start/$entry
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/ptr_deref_941_Split/split_ack
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/ptr_deref_941_Split/split_req
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/ptr_deref_941_Split/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/ptr_deref_941_Split/$entry
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/$entry
      -- 
    rr_2329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(214), ack => ptr_deref_941_store_0_req_0); -- 
    testConfigure_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(181) & testConfigure_CP_0_elements(185) & testConfigure_CP_0_elements(189) & testConfigure_CP_0_elements(193) & testConfigure_CP_0_elements(197) & testConfigure_CP_0_elements(201) & testConfigure_CP_0_elements(205) & testConfigure_CP_0_elements(209) & testConfigure_CP_0_elements(213);
      gj_testConfigure_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (5) 
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/word_access_start/word_0/ra
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/word_access_start/word_0/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/word_access_start/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Sample/$exit
      -- 
    ra_2330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_941_store_0_ack_0, ack => testConfigure_CP_0_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	289 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (5) 
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Update/word_access_complete/word_0/ca
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Update/word_access_complete/word_0/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Update/word_access_complete/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Update/$exit
      -- 
    ca_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_941_store_0_ack_1, ack => testConfigure_CP_0_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	178 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954__exit__
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_955__entry__
      -- CP-element group 217: 	 branch_block_stmt_32/R_exitcond8_956_place
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_955_else_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_955_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_955_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_955_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_955_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/if_stmt_955_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/$exit
      -- 
    branch_req_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(217), ack => if_stmt_955_branch_req_0); -- 
    testConfigure_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(178) & testConfigure_CP_0_elements(216);
      gj_testConfigure_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  transition  place  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	290 
    -- CP-element group 218:  members (13) 
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_961__exit__
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend189x_xloopexit_forx_xend189
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xbody135_forx_xend189x_xloopexit
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_955_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_955_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xbody135_forx_xend189x_xloopexit_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xbody135_forx_xend189x_xloopexit_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_961_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_961_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_961_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/merge_stmt_961_PhiAck/dummy
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend189x_xloopexit_forx_xend189_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/forx_xend189x_xloopexit_forx_xend189_PhiReq/$exit
      -- 
    if_choice_transition_2354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_955_branch_ack_1, ack => testConfigure_CP_0_elements(218)); -- 
    -- CP-element group 219:  fork  transition  place  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	285 
    -- CP-element group 219: 	286 
    -- CP-element group 219:  members (12) 
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_955_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_955_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/Sample/rr
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_955_branch_ack_0, ack => testConfigure_CP_0_elements(219)); -- 
    rr_2890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_798_inst_req_0); -- 
    cr_2895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_798_inst_req_1); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	290 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_Sample/ra
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_sample_completed_
      -- 
    ra_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_966_inst_ack_0, ack => testConfigure_CP_0_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	290 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (16) 
      -- CP-element group 221: 	 $exit
      -- CP-element group 221: 	 branch_block_stmt_32/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_967__exit__
      -- CP-element group 221: 	 branch_block_stmt_32/return__
      -- CP-element group 221: 	 branch_block_stmt_32/merge_stmt_969__exit__
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_967/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/merge_stmt_969_PhiReqMerge
      -- CP-element group 221: 	 branch_block_stmt_32/merge_stmt_969_PhiAck/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/merge_stmt_969_PhiAck/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/merge_stmt_969_PhiAck/dummy
      -- 
    ca_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_966_inst_ack_1, ack => testConfigure_CP_0_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	34 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (2) 
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/ra
      -- 
    ra_2409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => testConfigure_CP_0_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	34 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (2) 
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/ca
      -- 
    ca_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => testConfigure_CP_0_elements(223)); -- 
    -- CP-element group 224:  join  transition  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	228 
    -- CP-element group 224:  members (5) 
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_req
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/$exit
      -- 
    phi_stmt_73_req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(224), ack => phi_stmt_73_req_0); -- 
    testConfigure_cp_element_group_224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(222) & testConfigure_CP_0_elements(223);
      gj_testConfigure_cp_element_group_224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	34 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/ra
      -- 
    ra_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_0, ack => testConfigure_CP_0_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	34 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/ca
      -- 
    ca_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_1, ack => testConfigure_CP_0_elements(226)); -- 
    -- CP-element group 227:  join  transition  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_req
      -- 
    phi_stmt_80_req_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_80_req_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(227), ack => phi_stmt_80_req_0); -- 
    testConfigure_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(225) & testConfigure_CP_0_elements(226);
      gj_testConfigure_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  join  transition  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	224 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	234 
    -- CP-element group 228:  members (1) 
      -- CP-element group 228: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(224) & testConfigure_CP_0_elements(227);
      gj_testConfigure_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  transition  output  delay-element  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	14 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	233 
    -- CP-element group 229:  members (4) 
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_79_konst_delay_trans
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_req
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/$exit
      -- 
    phi_stmt_73_req_2449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_req_2449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => phi_stmt_73_req_1); -- 
    -- Element group testConfigure_CP_0_elements(229) is a control-delay.
    cp_element_229_delay: control_delay_element  generic map(name => " 229_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(14), ack => testConfigure_CP_0_elements(229), clk => clk, reset =>reset);
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	14 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (2) 
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/ra
      -- 
    ra_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_0, ack => testConfigure_CP_0_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	14 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (2) 
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/ca
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/$exit
      -- 
    ca_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_1, ack => testConfigure_CP_0_elements(231)); -- 
    -- CP-element group 232:  join  transition  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (5) 
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_req
      -- 
    phi_stmt_80_req_2472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_80_req_2472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(232), ack => phi_stmt_80_req_1); -- 
    testConfigure_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(230) & testConfigure_CP_0_elements(231);
      gj_testConfigure_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  transition  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	229 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(229) & testConfigure_CP_0_elements(232);
      gj_testConfigure_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  merge  fork  transition  place  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	228 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_32/merge_stmt_72_PhiReqMerge
      -- CP-element group 234: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(234) <= OrReduce(testConfigure_CP_0_elements(228) & testConfigure_CP_0_elements(233));
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (1) 
      -- CP-element group 235: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/phi_stmt_73_ack
      -- 
    phi_stmt_73_ack_2477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_73_ack_0, ack => testConfigure_CP_0_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/phi_stmt_80_ack
      -- 
    phi_stmt_80_ack_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_80_ack_0, ack => testConfigure_CP_0_elements(236)); -- 
    -- CP-element group 237:  join  fork  transition  place  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	15 
    -- CP-element group 237: 	16 
    -- CP-element group 237: 	17 
    -- CP-element group 237: 	18 
    -- CP-element group 237: 	20 
    -- CP-element group 237: 	22 
    -- CP-element group 237: 	23 
    -- CP-element group 237: 	25 
    -- CP-element group 237: 	27 
    -- CP-element group 237: 	28 
    -- CP-element group 237: 	31 
    -- CP-element group 237:  members (64) 
      -- CP-element group 237: 	 branch_block_stmt_32/merge_stmt_72__exit__
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142__entry__
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_addrgen/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_addrgen/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_addrgen/root_register_req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_addrgen/root_register_ack
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Sample/rr
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_95_Update/cr
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resized_1
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scaled_1
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_computed_1
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resize_1/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resize_1/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resize_1/index_resize_req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_resize_1/index_resize_ack
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scale_1/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scale_1/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scale_1/scale_rename_req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_index_scale_1/scale_rename_ack
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_update_start
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Sample/req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/array_obj_ref_101_final_index_sum_regn_Update/req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_complete/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/addr_of_102_complete/req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/word_0/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_105_Update/word_access_complete/word_0/cr
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_address_calculated
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_word_address_calculated
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_root_address_calculated
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_address_resized
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_addr_resize/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_addr_resize/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_addr_resize/base_resize_req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_addr_resize/base_resize_ack
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_plus_offset/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_plus_offset/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_plus_offset/sum_rename_req
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_base_plus_offset/sum_rename_ack
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/word_0/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/ptr_deref_122_Update/word_access_complete/word_0/cr
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_126_Update/cr
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/RPIPE_ConvTranspose_input_pipe_137_Sample/rr
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_142/type_cast_141_Update/cr
      -- CP-element group 237: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/$exit
      -- 
    rr_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => type_cast_95_inst_req_0); -- 
    cr_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => type_cast_95_inst_req_1); -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => array_obj_ref_101_index_offset_req_0); -- 
    req_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => array_obj_ref_101_index_offset_req_1); -- 
    req_279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => addr_of_102_final_reg_req_1); -- 
    cr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => ptr_deref_105_store_0_req_1); -- 
    cr_374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => ptr_deref_122_load_0_req_1); -- 
    cr_393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => type_cast_126_inst_req_1); -- 
    rr_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => RPIPE_ConvTranspose_input_pipe_137_inst_req_0); -- 
    cr_421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(237), ack => type_cast_141_inst_req_1); -- 
    testConfigure_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(235) & testConfigure_CP_0_elements(236);
      gj_testConfigure_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	35 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (2) 
      -- CP-element group 238: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/ra
      -- CP-element group 238: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/$exit
      -- 
    ra_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_0, ack => testConfigure_CP_0_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	35 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/ca
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/$exit
      -- 
    ca_2507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_1, ack => testConfigure_CP_0_elements(239)); -- 
    -- CP-element group 240:  join  transition  place  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (8) 
      -- CP-element group 240: 	 branch_block_stmt_32/merge_stmt_149_PhiReqMerge
      -- CP-element group 240: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/$entry
      -- CP-element group 240: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_req
      -- CP-element group 240: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/phi_stmt_150_sources/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_150/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- 
    phi_stmt_150_req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(240), ack => phi_stmt_150_req_0); -- 
    testConfigure_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(238) & testConfigure_CP_0_elements(239);
      gj_testConfigure_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	245 
    -- CP-element group 241: 	246 
    -- CP-element group 241:  members (13) 
      -- CP-element group 241: 	 branch_block_stmt_32/merge_stmt_149__exit__
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Update/cr
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Sample/rr
      -- CP-element group 241: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/phi_stmt_150_ack
      -- CP-element group 241: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/$entry
      -- 
    phi_stmt_150_ack_2513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_150_ack_0, ack => testConfigure_CP_0_elements(241)); -- 
    cr_2563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => type_cast_162_inst_req_1); -- 
    rr_2558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => type_cast_162_inst_req_0); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	13 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Sample/ra
      -- CP-element group 242: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Sample/$exit
      -- 
    ra_2533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_160_inst_ack_0, ack => testConfigure_CP_0_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	13 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/Update/ca
      -- 
    ca_2538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_160_inst_ack_1, ack => testConfigure_CP_0_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	248 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_req
      -- CP-element group 244: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/SplitProtocol/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_160/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_157/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_157_req_2539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_157_req_2539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => phi_stmt_157_req_0); -- 
    testConfigure_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(242) & testConfigure_CP_0_elements(243);
      gj_testConfigure_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	241 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (2) 
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Sample/ra
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Sample/$exit
      -- 
    ra_2559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_162_inst_ack_0, ack => testConfigure_CP_0_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	241 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Update/ca
      -- CP-element group 246: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/Update/$exit
      -- 
    ca_2564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_162_inst_ack_1, ack => testConfigure_CP_0_elements(246)); -- 
    -- CP-element group 247:  join  transition  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_req
      -- CP-element group 247: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/SplitProtocol/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/type_cast_162/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/phi_stmt_157_sources/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_157/$exit
      -- 
    phi_stmt_157_req_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_157_req_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(247), ack => phi_stmt_157_req_1); -- 
    testConfigure_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(245) & testConfigure_CP_0_elements(246);
      gj_testConfigure_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  merge  transition  place  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	244 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (2) 
      -- CP-element group 248: 	 branch_block_stmt_32/merge_stmt_156_PhiReqMerge
      -- CP-element group 248: 	 branch_block_stmt_32/merge_stmt_156_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(248) <= OrReduce(testConfigure_CP_0_elements(244) & testConfigure_CP_0_elements(247));
    -- CP-element group 249:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	36 
    -- CP-element group 249: 	37 
    -- CP-element group 249:  members (35) 
      -- CP-element group 249: 	 branch_block_stmt_32/merge_stmt_156__exit__
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179__entry__
      -- CP-element group 249: 	 branch_block_stmt_32/merge_stmt_156_PhiAck/phi_stmt_157_ack
      -- CP-element group 249: 	 branch_block_stmt_32/merge_stmt_156_PhiAck/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_root_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_address_resized
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_addr_resize/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_addr_resize/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_addr_resize/base_resize_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_addr_resize/base_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_plus_offset/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_plus_offset/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_plus_offset/sum_rename_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_base_plus_offset/sum_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_addrgen/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_addrgen/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_addrgen/root_register_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_word_addrgen/root_register_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/ptr_deref_171_Split/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/ptr_deref_171_Split/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/ptr_deref_171_Split/split_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/ptr_deref_171_Split/split_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Sample/word_access_start/word_0/rr
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_169_to_assign_stmt_179/ptr_deref_171_Update/word_access_complete/word_0/cr
      -- 
    phi_stmt_157_ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_157_ack_0, ack => testConfigure_CP_0_elements(249)); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => ptr_deref_171_store_0_req_0); -- 
    cr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => ptr_deref_171_store_0_req_1); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	60 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Sample/ra
      -- CP-element group 250: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Sample/$exit
      -- 
    ra_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_0, ack => testConfigure_CP_0_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	60 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Update/ca
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/Update/$exit
      -- 
    ca_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_192_inst_ack_1, ack => testConfigure_CP_0_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_req
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_192/SplitProtocol/$exit
      -- 
    phi_stmt_189_req_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_189_req_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(252), ack => phi_stmt_189_req_0); -- 
    testConfigure_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(250) & testConfigure_CP_0_elements(251);
      gj_testConfigure_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  transition  output  delay-element  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	39 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (5) 
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_req
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_189/phi_stmt_189_sources/type_cast_195_konst_delay_trans
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/$exit
      -- 
    phi_stmt_189_req_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_189_req_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => phi_stmt_189_req_1); -- 
    -- Element group testConfigure_CP_0_elements(253) is a control-delay.
    cp_element_253_delay: control_delay_element  generic map(name => " 253_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(39), ack => testConfigure_CP_0_elements(253), clk => clk, reset =>reset);
    -- CP-element group 254:  merge  transition  place  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_32/merge_stmt_188_PhiReqMerge
      -- CP-element group 254: 	 branch_block_stmt_32/merge_stmt_188_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(254) <= OrReduce(testConfigure_CP_0_elements(252) & testConfigure_CP_0_elements(253));
    -- CP-element group 255:  fork  transition  place  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	40 
    -- CP-element group 255: 	41 
    -- CP-element group 255: 	42 
    -- CP-element group 255: 	43 
    -- CP-element group 255: 	45 
    -- CP-element group 255: 	46 
    -- CP-element group 255: 	49 
    -- CP-element group 255: 	52 
    -- CP-element group 255: 	53 
    -- CP-element group 255: 	55 
    -- CP-element group 255: 	57 
    -- CP-element group 255:  members (65) 
      -- CP-element group 255: 	 branch_block_stmt_32/merge_stmt_188__exit__
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251__entry__
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Sample/rr
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_205_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resized_1
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scaled_1
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_computed_1
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resize_1/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resize_1/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resize_1/index_resize_req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_resize_1/index_resize_ack
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scale_1/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scale_1/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scale_1/scale_rename_req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_index_scale_1/scale_rename_ack
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_update_start
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Sample/req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/array_obj_ref_211_final_index_sum_regn_Update/req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_complete/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/addr_of_212_complete/req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/RPIPE_ConvTranspose_input_pipe_215_Sample/rr
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_219_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/word_0/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_222_Update/word_access_complete/word_0/cr
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_address_calculated
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_address_calculated
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_root_address_calculated
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_address_resized
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_addr_resize/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_addr_resize/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_addr_resize/base_resize_req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_addr_resize/base_resize_ack
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_plus_offset/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_plus_offset/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_plus_offset/sum_rename_req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_base_plus_offset/sum_rename_ack
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_addrgen/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_addrgen/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_addrgen/root_register_req
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_word_addrgen/root_register_ack
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/word_0/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/ptr_deref_239_Update/word_access_complete/word_0/cr
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/assign_stmt_202_to_assign_stmt_251/type_cast_243_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_32/merge_stmt_188_PhiAck/phi_stmt_189_ack
      -- CP-element group 255: 	 branch_block_stmt_32/merge_stmt_188_PhiAck/$exit
      -- 
    phi_stmt_189_ack_2624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_189_ack_0, ack => testConfigure_CP_0_elements(255)); -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => type_cast_205_inst_req_0); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => type_cast_205_inst_req_1); -- 
    req_556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => array_obj_ref_211_index_offset_req_0); -- 
    req_561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => array_obj_ref_211_index_offset_req_1); -- 
    req_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => addr_of_212_final_reg_req_1); -- 
    rr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => RPIPE_ConvTranspose_input_pipe_215_inst_req_0); -- 
    cr_604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => type_cast_219_inst_req_1); -- 
    cr_654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => ptr_deref_222_store_0_req_1); -- 
    cr_699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => ptr_deref_239_load_0_req_1); -- 
    cr_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => type_cast_243_inst_req_1); -- 
    -- CP-element group 256:  merge  fork  transition  place  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	38 
    -- CP-element group 256: 	61 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	62 
    -- CP-element group 256: 	65 
    -- CP-element group 256:  members (13) 
      -- CP-element group 256: 	 branch_block_stmt_32/merge_stmt_260__exit__
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267__entry__
      -- CP-element group 256: 	 branch_block_stmt_32/merge_stmt_260_PhiAck/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/merge_stmt_260_PhiAck/dummy
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/RPIPE_ConvTranspose_input_pipe_262_Sample/rr
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_update_start_
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/assign_stmt_263_to_assign_stmt_267/type_cast_266_Update/cr
      -- CP-element group 256: 	 branch_block_stmt_32/merge_stmt_260_PhiReqMerge
      -- CP-element group 256: 	 branch_block_stmt_32/merge_stmt_260_PhiAck/$entry
      -- 
    rr_750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(256), ack => RPIPE_ConvTranspose_input_pipe_262_inst_req_0); -- 
    cr_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(256), ack => type_cast_266_inst_req_1); -- 
    testConfigure_CP_0_elements(256) <= OrReduce(testConfigure_CP_0_elements(38) & testConfigure_CP_0_elements(61));
    -- CP-element group 257:  transition  output  delay-element  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	65 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	261 
    -- CP-element group 257:  members (4) 
      -- CP-element group 257: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_270/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_274_konst_delay_trans
      -- CP-element group 257: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_req
      -- 
    phi_stmt_270_req_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_270_req_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(257), ack => phi_stmt_270_req_0); -- 
    -- Element group testConfigure_CP_0_elements(257) is a control-delay.
    cp_element_257_delay: control_delay_element  generic map(name => " 257_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(65), ack => testConfigure_CP_0_elements(257), clk => clk, reset =>reset);
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	65 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Sample/ra
      -- 
    ra_2675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_0, ack => testConfigure_CP_0_elements(258)); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	65 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (2) 
      -- CP-element group 259: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/Update/ca
      -- 
    ca_2680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_1, ack => testConfigure_CP_0_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (5) 
      -- CP-element group 260: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_280/SplitProtocol/$exit
      -- CP-element group 260: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_req
      -- 
    phi_stmt_277_req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_277_req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(260), ack => phi_stmt_277_req_0); -- 
    testConfigure_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(258) & testConfigure_CP_0_elements(259);
      gj_testConfigure_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  join  transition  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	257 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	269 
    -- CP-element group 261:  members (1) 
      -- CP-element group 261: 	 branch_block_stmt_32/bbx_xnph207_forx_xbody30_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(257) & testConfigure_CP_0_elements(260);
      gj_testConfigure_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	76 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (2) 
      -- CP-element group 262: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Sample/ra
      -- 
    ra_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_276_inst_ack_0, ack => testConfigure_CP_0_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	76 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (2) 
      -- CP-element group 263: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/Update/ca
      -- 
    ca_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_276_inst_ack_1, ack => testConfigure_CP_0_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	268 
    -- CP-element group 264:  members (5) 
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_sources/type_cast_276/SplitProtocol/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_270/phi_stmt_270_req
      -- 
    phi_stmt_270_req_2707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_270_req_2707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => phi_stmt_270_req_1); -- 
    testConfigure_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(262) & testConfigure_CP_0_elements(263);
      gj_testConfigure_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	76 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (2) 
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Sample/ra
      -- 
    ra_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_282_inst_ack_0, ack => testConfigure_CP_0_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	76 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/Update/ca
      -- 
    ca_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_282_inst_ack_1, ack => testConfigure_CP_0_elements(266)); -- 
    -- CP-element group 267:  join  transition  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (5) 
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_sources/type_cast_282/SplitProtocol/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/phi_stmt_277/phi_stmt_277_req
      -- 
    phi_stmt_277_req_2730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_277_req_2730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => phi_stmt_277_req_1); -- 
    testConfigure_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(265) & testConfigure_CP_0_elements(266);
      gj_testConfigure_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  join  transition  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	264 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (1) 
      -- CP-element group 268: 	 branch_block_stmt_32/forx_xbody30_forx_xbody30_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(264) & testConfigure_CP_0_elements(267);
      gj_testConfigure_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  merge  fork  transition  place  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	261 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (2) 
      -- CP-element group 269: 	 branch_block_stmt_32/merge_stmt_269_PhiReqMerge
      -- CP-element group 269: 	 branch_block_stmt_32/merge_stmt_269_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(269) <= OrReduce(testConfigure_CP_0_elements(261) & testConfigure_CP_0_elements(268));
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (1) 
      -- CP-element group 270: 	 branch_block_stmt_32/merge_stmt_269_PhiAck/phi_stmt_270_ack
      -- 
    phi_stmt_270_ack_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_270_ack_0, ack => testConfigure_CP_0_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (1) 
      -- CP-element group 271: 	 branch_block_stmt_32/merge_stmt_269_PhiAck/phi_stmt_277_ack
      -- 
    phi_stmt_277_ack_2736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_277_ack_0, ack => testConfigure_CP_0_elements(271)); -- 
    -- CP-element group 272:  join  fork  transition  place  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	66 
    -- CP-element group 272: 	67 
    -- CP-element group 272: 	69 
    -- CP-element group 272: 	70 
    -- CP-element group 272: 	73 
    -- CP-element group 272:  members (42) 
      -- CP-element group 272: 	 branch_block_stmt_32/merge_stmt_269__exit__
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311__entry__
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scale_0/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scale_0/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scale_0/scale_rename_req
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scale_0/scale_rename_ack
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_final_index_sum_regn/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_final_index_sum_regn/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_final_index_sum_regn/req
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_final_index_sum_regn/ack
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_base_plus_offset/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_base_plus_offset/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_base_plus_offset/sum_rename_req
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_base_plus_offset/sum_rename_ack
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_request/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_request/req
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_complete/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_complete/req
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/addr_of_287_update_start_
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_root_address_calculated
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_offset_calculated
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resized_0
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_scaled_0
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_computed_0
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resize_0/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resize_0/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resize_0/index_resize_req
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/array_obj_ref_286_index_resize_0/index_resize_ack
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_update_start_
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/word_0/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/ptr_deref_290_Update/word_access_complete/word_0/cr
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/RPIPE_ConvTranspose_input_pipe_294_Sample/rr
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_update_start_
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/assign_stmt_288_to_assign_stmt_311/type_cast_298_Update/cr
      -- CP-element group 272: 	 branch_block_stmt_32/merge_stmt_269_PhiAck/$exit
      -- 
    req_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => addr_of_287_final_reg_req_0); -- 
    req_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => addr_of_287_final_reg_req_1); -- 
    cr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => ptr_deref_290_store_0_req_1); -- 
    rr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => RPIPE_ConvTranspose_input_pipe_294_inst_req_0); -- 
    cr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => type_cast_298_inst_req_1); -- 
    testConfigure_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(270) & testConfigure_CP_0_elements(271);
      gj_testConfigure_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	75 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (2) 
      -- CP-element group 273: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Sample/ra
      -- 
    ra_2760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_0, ack => testConfigure_CP_0_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	75 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/Update/ca
      -- 
    ca_2765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_1, ack => testConfigure_CP_0_elements(274)); -- 
    -- CP-element group 275:  join  transition  place  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (8) 
      -- CP-element group 275: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_sources/type_cast_322/SplitProtocol/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/forx_xbody30_forx_xend39_PhiReq/phi_stmt_319/phi_stmt_319_req
      -- CP-element group 275: 	 branch_block_stmt_32/merge_stmt_318_PhiReqMerge
      -- CP-element group 275: 	 branch_block_stmt_32/merge_stmt_318_PhiAck/$entry
      -- 
    phi_stmt_319_req_2766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_319_req_2766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => phi_stmt_319_req_0); -- 
    testConfigure_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(273) & testConfigure_CP_0_elements(274);
      gj_testConfigure_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  merge  transition  place  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	77 
    -- CP-element group 276:  members (4) 
      -- CP-element group 276: 	 branch_block_stmt_32/merge_stmt_318__exit__
      -- CP-element group 276: 	 branch_block_stmt_32/assign_stmt_326_to_assign_stmt_557__entry__
      -- CP-element group 276: 	 branch_block_stmt_32/merge_stmt_318_PhiAck/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/merge_stmt_318_PhiAck/phi_stmt_319_ack
      -- 
    phi_stmt_319_ack_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_319_ack_0, ack => testConfigure_CP_0_elements(276)); -- 
    -- CP-element group 277:  merge  branch  transition  place  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	133 
    -- CP-element group 277: 	176 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	134 
    -- CP-element group 277: 	135 
    -- CP-element group 277:  members (17) 
      -- CP-element group 277: 	 branch_block_stmt_32/merge_stmt_566__exit__
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_572__entry__
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_572__exit__
      -- CP-element group 277: 	 branch_block_stmt_32/if_stmt_573__entry__
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_572/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/assign_stmt_572/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/if_stmt_573_dead_link/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/if_stmt_573_eval_test/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/if_stmt_573_eval_test/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/if_stmt_573_eval_test/branch_req
      -- CP-element group 277: 	 branch_block_stmt_32/R_cmp133195_574_place
      -- CP-element group 277: 	 branch_block_stmt_32/if_stmt_573_if_link/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/if_stmt_573_else_link/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/merge_stmt_566_PhiReqMerge
      -- CP-element group 277: 	 branch_block_stmt_32/merge_stmt_566_PhiAck/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/merge_stmt_566_PhiAck/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/merge_stmt_566_PhiAck/dummy
      -- 
    branch_req_1659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => if_stmt_573_branch_req_0); -- 
    testConfigure_CP_0_elements(277) <= OrReduce(testConfigure_CP_0_elements(133) & testConfigure_CP_0_elements(176));
    -- CP-element group 278:  transition  output  delay-element  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	132 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	282 
    -- CP-element group 278:  members (5) 
      -- CP-element group 278: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76_PhiReq/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76_PhiReq/phi_stmt_601/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_605_konst_delay_trans
      -- CP-element group 278: 	 branch_block_stmt_32/bbx_xnph201_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_req
      -- 
    phi_stmt_601_req_2817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_601_req_2817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(278), ack => phi_stmt_601_req_0); -- 
    -- Element group testConfigure_CP_0_elements(278) is a control-delay.
    cp_element_278_delay: control_delay_element  generic map(name => " 278_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(132), ack => testConfigure_CP_0_elements(278), clk => clk, reset =>reset);
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	177 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (2) 
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/Sample/ra
      -- 
    ra_2837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_607_inst_ack_0, ack => testConfigure_CP_0_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	177 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (2) 
      -- CP-element group 280: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/Update/ca
      -- 
    ca_2842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_607_inst_ack_1, ack => testConfigure_CP_0_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_sources/type_cast_607/SplitProtocol/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/forx_xbody76_forx_xbody76_PhiReq/phi_stmt_601/phi_stmt_601_req
      -- 
    phi_stmt_601_req_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_601_req_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(281), ack => phi_stmt_601_req_1); -- 
    testConfigure_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(279) & testConfigure_CP_0_elements(280);
      gj_testConfigure_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  merge  transition  place  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	278 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (2) 
      -- CP-element group 282: 	 branch_block_stmt_32/merge_stmt_600_PhiReqMerge
      -- CP-element group 282: 	 branch_block_stmt_32/merge_stmt_600_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(282) <= OrReduce(testConfigure_CP_0_elements(278) & testConfigure_CP_0_elements(281));
    -- CP-element group 283:  fork  transition  place  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	136 
    -- CP-element group 283: 	137 
    -- CP-element group 283: 	139 
    -- CP-element group 283: 	140 
    -- CP-element group 283: 	143 
    -- CP-element group 283: 	147 
    -- CP-element group 283: 	151 
    -- CP-element group 283: 	155 
    -- CP-element group 283: 	159 
    -- CP-element group 283: 	163 
    -- CP-element group 283: 	167 
    -- CP-element group 283: 	171 
    -- CP-element group 283: 	174 
    -- CP-element group 283:  members (56) 
      -- CP-element group 283: 	 branch_block_stmt_32/merge_stmt_600__exit__
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763__entry__
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_resized_1
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_scaled_1
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_computed_1
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_resize_1/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_resize_1/$exit
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_resize_1/index_resize_req
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_resize_1/index_resize_ack
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_scale_1/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_scale_1/$exit
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_scale_1/scale_rename_req
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_index_scale_1/scale_rename_ack
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_update_start
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/array_obj_ref_613_final_index_sum_regn_Update/req
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_complete/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/addr_of_614_complete/req
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/RPIPE_ConvTranspose_input_pipe_617_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_621_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_634_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_652_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_670_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_688_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_706_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_724_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/type_cast_742_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Update/word_access_complete/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Update/word_access_complete/word_0/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/assign_stmt_615_to_assign_stmt_763/ptr_deref_750_Update/word_access_complete/word_0/cr
      -- CP-element group 283: 	 branch_block_stmt_32/merge_stmt_600_PhiAck/$exit
      -- CP-element group 283: 	 branch_block_stmt_32/merge_stmt_600_PhiAck/phi_stmt_601_ack
      -- 
    phi_stmt_601_ack_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_601_ack_0, ack => testConfigure_CP_0_elements(283)); -- 
    req_1701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => array_obj_ref_613_index_offset_req_0); -- 
    req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => array_obj_ref_613_index_offset_req_1); -- 
    req_1721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => addr_of_614_final_reg_req_1); -- 
    rr_1730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => RPIPE_ConvTranspose_input_pipe_617_inst_req_0); -- 
    cr_1749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_621_inst_req_1); -- 
    cr_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_634_inst_req_1); -- 
    cr_1805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_652_inst_req_1); -- 
    cr_1833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_670_inst_req_1); -- 
    cr_1861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_688_inst_req_1); -- 
    cr_1889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_706_inst_req_1); -- 
    cr_1917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_724_inst_req_1); -- 
    cr_1945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => type_cast_742_inst_req_1); -- 
    cr_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => ptr_deref_750_store_0_req_1); -- 
    -- CP-element group 284:  transition  output  delay-element  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	134 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	288 
    -- CP-element group 284:  members (5) 
      -- CP-element group 284: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135_PhiReq/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135_PhiReq/phi_stmt_792/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_796_konst_delay_trans
      -- CP-element group 284: 	 branch_block_stmt_32/bbx_xnph_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_req
      -- 
    phi_stmt_792_req_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_792_req_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => phi_stmt_792_req_0); -- 
    -- Element group testConfigure_CP_0_elements(284) is a control-delay.
    cp_element_284_delay: control_delay_element  generic map(name => " 284_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(134), ack => testConfigure_CP_0_elements(284), clk => clk, reset =>reset);
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	219 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/Sample/ra
      -- 
    ra_2891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_798_inst_ack_0, ack => testConfigure_CP_0_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	219 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/Update/ca
      -- 
    ca_2896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_798_inst_ack_1, ack => testConfigure_CP_0_elements(286)); -- 
    -- CP-element group 287:  join  transition  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (6) 
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_sources/type_cast_798/SplitProtocol/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody135_forx_xbody135_PhiReq/phi_stmt_792/phi_stmt_792_req
      -- 
    phi_stmt_792_req_2897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_792_req_2897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => phi_stmt_792_req_1); -- 
    testConfigure_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(285) & testConfigure_CP_0_elements(286);
      gj_testConfigure_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  merge  transition  place  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	284 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (2) 
      -- CP-element group 288: 	 branch_block_stmt_32/merge_stmt_791_PhiReqMerge
      -- CP-element group 288: 	 branch_block_stmt_32/merge_stmt_791_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(288) <= OrReduce(testConfigure_CP_0_elements(284) & testConfigure_CP_0_elements(287));
    -- CP-element group 289:  fork  transition  place  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	178 
    -- CP-element group 289: 	179 
    -- CP-element group 289: 	181 
    -- CP-element group 289: 	182 
    -- CP-element group 289: 	185 
    -- CP-element group 289: 	189 
    -- CP-element group 289: 	193 
    -- CP-element group 289: 	197 
    -- CP-element group 289: 	201 
    -- CP-element group 289: 	205 
    -- CP-element group 289: 	209 
    -- CP-element group 289: 	213 
    -- CP-element group 289: 	216 
    -- CP-element group 289:  members (56) 
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_32/merge_stmt_791__exit__
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954__entry__
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_933_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_879_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_915_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Update/word_access_complete/word_0/cr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Update/word_access_complete/word_0/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Update/word_access_complete/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/ptr_deref_941_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_897_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_resized_1
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_scaled_1
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_computed_1
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_resize_1/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_resize_1/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_resize_1/index_resize_req
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_resize_1/index_resize_ack
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_scale_1/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_scale_1/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_scale_1/scale_rename_req
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_index_scale_1/scale_rename_ack
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_update_start
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_Sample/req
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/array_obj_ref_804_final_index_sum_regn_Update/req
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_complete/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/addr_of_805_complete/req
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/RPIPE_ConvTranspose_input_pipe_808_Sample/rr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_812_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_825_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_843_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_806_to_assign_stmt_954/type_cast_861_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/merge_stmt_791_PhiAck/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/merge_stmt_791_PhiAck/phi_stmt_792_ack
      -- 
    phi_stmt_792_ack_2902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_792_ack_0, ack => testConfigure_CP_0_elements(289)); -- 
    cr_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => type_cast_861_inst_req_1); -- 
    cr_2262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => type_cast_915_inst_req_1); -- 
    cr_2290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => type_cast_933_inst_req_1); -- 
    cr_2206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => type_cast_879_inst_req_1); -- 
    cr_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => ptr_deref_941_store_0_req_1); -- 
    cr_2234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => type_cast_897_inst_req_1); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => array_obj_ref_804_index_offset_req_0); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => array_obj_ref_804_index_offset_req_1); -- 
    req_2066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => addr_of_805_final_reg_req_1); -- 
    rr_2075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => RPIPE_ConvTranspose_input_pipe_808_inst_req_0); -- 
    cr_2094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => type_cast_812_inst_req_1); -- 
    cr_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => type_cast_825_inst_req_1); -- 
    cr_2150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => type_cast_843_inst_req_1); -- 
    -- CP-element group 290:  merge  fork  transition  place  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	135 
    -- CP-element group 290: 	218 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	220 
    -- CP-element group 290: 	221 
    -- CP-element group 290:  members (13) 
      -- CP-element group 290: 	 branch_block_stmt_32/merge_stmt_963__exit__
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_967__entry__
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_Sample/rr
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_update_start_
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_967/type_cast_966_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_32/assign_stmt_967/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/merge_stmt_963_PhiReqMerge
      -- CP-element group 290: 	 branch_block_stmt_32/merge_stmt_963_PhiAck/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/merge_stmt_963_PhiAck/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/merge_stmt_963_PhiAck/dummy
      -- 
    cr_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(290), ack => type_cast_966_inst_req_1); -- 
    rr_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(290), ack => type_cast_966_inst_req_0); -- 
    testConfigure_CP_0_elements(290) <= OrReduce(testConfigure_CP_0_elements(135) & testConfigure_CP_0_elements(218));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_455_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_549_wire : std_logic_vector(63 downto 0);
    signal R_indvar222_612_resized : std_logic_vector(13 downto 0);
    signal R_indvar222_612_scaled : std_logic_vector(13 downto 0);
    signal R_indvar228_285_resized : std_logic_vector(0 downto 0);
    signal R_indvar228_285_scaled : std_logic_vector(0 downto 0);
    signal R_indvar231_210_resized : std_logic_vector(6 downto 0);
    signal R_indvar231_210_scaled : std_logic_vector(6 downto 0);
    signal R_indvar236_100_resized : std_logic_vector(6 downto 0);
    signal R_indvar236_100_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_803_resized : std_logic_vector(10 downto 0);
    signal R_indvar_803_scaled : std_logic_vector(10 downto 0);
    signal STORE_padding_324_data_0 : std_logic_vector(15 downto 0);
    signal STORE_padding_324_word_address_0 : std_logic_vector(0 downto 0);
    signal add101_694 : std_logic_vector(63 downto 0);
    signal add107_712 : std_logic_vector(63 downto 0);
    signal add113_730 : std_logic_vector(63 downto 0);
    signal add119_748 : std_logic_vector(63 downto 0);
    signal add145_831 : std_logic_vector(63 downto 0);
    signal add151_849 : std_logic_vector(63 downto 0);
    signal add157_867 : std_logic_vector(63 downto 0);
    signal add163_885 : std_logic_vector(63 downto 0);
    signal add169_903 : std_logic_vector(63 downto 0);
    signal add175_921 : std_logic_vector(63 downto 0);
    signal add181_939 : std_logic_vector(63 downto 0);
    signal add89_658 : std_logic_vector(63 downto 0);
    signal add95_676 : std_logic_vector(63 downto 0);
    signal add_640 : std_logic_vector(63 downto 0);
    signal array_obj_ref_101_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_211_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_286_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_286_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_286_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_286_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_613_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_613_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_613_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_613_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_613_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_613_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_804_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_804_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_804_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_804_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_804_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_804_root_address : std_logic_vector(10 downto 0);
    signal arrayidx123_615 : std_logic_vector(31 downto 0);
    signal arrayidx185_806 : std_logic_vector(31 downto 0);
    signal arrayidx21_213 : std_logic_vector(31 downto 0);
    signal arrayidx35_288 : std_logic_vector(31 downto 0);
    signal arrayidx_103 : std_logic_vector(31 downto 0);
    signal call104_703 : std_logic_vector(7 downto 0);
    signal call110_721 : std_logic_vector(7 downto 0);
    signal call116_739 : std_logic_vector(7 downto 0);
    signal call138_809 : std_logic_vector(7 downto 0);
    signal call142_822 : std_logic_vector(7 downto 0);
    signal call148_840 : std_logic_vector(7 downto 0);
    signal call154_858 : std_logic_vector(7 downto 0);
    signal call160_876 : std_logic_vector(7 downto 0);
    signal call166_894 : std_logic_vector(7 downto 0);
    signal call172_912 : std_logic_vector(7 downto 0);
    signal call178_930 : std_logic_vector(7 downto 0);
    signal call17_216 : std_logic_vector(7 downto 0);
    signal call31203_263 : std_logic_vector(7 downto 0);
    signal call31_295 : std_logic_vector(7 downto 0);
    signal call4216_59 : std_logic_vector(7 downto 0);
    signal call42_329 : std_logic_vector(7 downto 0);
    signal call44_348 : std_logic_vector(7 downto 0);
    signal call46_367 : std_logic_vector(7 downto 0);
    signal call4_138 : std_logic_vector(7 downto 0);
    signal call78_618 : std_logic_vector(7 downto 0);
    signal call81_631 : std_logic_vector(7 downto 0);
    signal call86_649 : std_logic_vector(7 downto 0);
    signal call92_667 : std_logic_vector(7 downto 0);
    signal call98_685 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp133195_572 : std_logic_vector(0 downto 0);
    signal cmp14210_179 : std_logic_vector(0 downto 0);
    signal cmp14_251 : std_logic_vector(0 downto 0);
    signal cmp215_56 : std_logic_vector(0 downto 0);
    signal cmp74199_557 : std_logic_vector(0 downto 0);
    signal cmp_135 : std_logic_vector(0 downto 0);
    signal conv100_689 : std_logic_vector(63 downto 0);
    signal conv106_707 : std_logic_vector(63 downto 0);
    signal conv112_725 : std_logic_vector(63 downto 0);
    signal conv118_743 : std_logic_vector(63 downto 0);
    signal conv139_813 : std_logic_vector(63 downto 0);
    signal conv13_244 : std_logic_vector(31 downto 0);
    signal conv144_826 : std_logic_vector(63 downto 0);
    signal conv150_844 : std_logic_vector(63 downto 0);
    signal conv156_862 : std_logic_vector(63 downto 0);
    signal conv162_880 : std_logic_vector(63 downto 0);
    signal conv168_898 : std_logic_vector(63 downto 0);
    signal conv174_916 : std_logic_vector(63 downto 0);
    signal conv180_934 : std_logic_vector(63 downto 0);
    signal conv18_220 : std_logic_vector(15 downto 0);
    signal conv2_127 : std_logic_vector(31 downto 0);
    signal conv32204_267 : std_logic_vector(15 downto 0);
    signal conv32206_277 : std_logic_vector(15 downto 0);
    signal conv32_299 : std_logic_vector(15 downto 0);
    signal conv32x_xlcssa_319 : std_logic_vector(15 downto 0);
    signal conv43_333 : std_logic_vector(15 downto 0);
    signal conv45_352 : std_logic_vector(15 downto 0);
    signal conv47_371 : std_logic_vector(15 downto 0);
    signal conv50_399 : std_logic_vector(63 downto 0);
    signal conv5217_63 : std_logic_vector(15 downto 0);
    signal conv5219_80 : std_logic_vector(15 downto 0);
    signal conv52_415 : std_logic_vector(63 downto 0);
    signal conv54_431 : std_logic_vector(63 downto 0);
    signal conv56_457 : std_logic_vector(63 downto 0);
    signal conv59_473 : std_logic_vector(63 downto 0);
    signal conv5_142 : std_logic_vector(15 downto 0);
    signal conv5x_xlcssa1_150 : std_logic_vector(15 downto 0);
    signal conv5x_xlcssa_157 : std_logic_vector(15 downto 0);
    signal conv61_489 : std_logic_vector(63 downto 0);
    signal conv64_505 : std_logic_vector(63 downto 0);
    signal conv67_521 : std_logic_vector(63 downto 0);
    signal conv69_551 : std_logic_vector(63 downto 0);
    signal conv79_622 : std_logic_vector(63 downto 0);
    signal conv83_635 : std_logic_vector(63 downto 0);
    signal conv88_653 : std_logic_vector(63 downto 0);
    signal conv94_671 : std_logic_vector(63 downto 0);
    signal conv_39 : std_logic_vector(15 downto 0);
    signal exitcond8_954 : std_logic_vector(0 downto 0);
    signal exitcond9_311 : std_logic_vector(0 downto 0);
    signal exitcond_763 : std_logic_vector(0 downto 0);
    signal iNsTr_13_119 : std_logic_vector(31 downto 0);
    signal iNsTr_1_45 : std_logic_vector(31 downto 0);
    signal iNsTr_21_236 : std_logic_vector(31 downto 0);
    signal iNsTr_26_341 : std_logic_vector(31 downto 0);
    signal iNsTr_29_360 : std_logic_vector(31 downto 0);
    signal iNsTr_32_379 : std_logic_vector(31 downto 0);
    signal iNsTr_34_391 : std_logic_vector(31 downto 0);
    signal iNsTr_35_407 : std_logic_vector(31 downto 0);
    signal iNsTr_36_423 : std_logic_vector(31 downto 0);
    signal iNsTr_37_465 : std_logic_vector(31 downto 0);
    signal iNsTr_38_481 : std_logic_vector(31 downto 0);
    signal iNsTr_39_497 : std_logic_vector(31 downto 0);
    signal iNsTr_40_513 : std_logic_vector(31 downto 0);
    signal iNsTr_5_169 : std_logic_vector(31 downto 0);
    signal inc24_206 : std_logic_vector(31 downto 0);
    signal inc_96 : std_logic_vector(31 downto 0);
    signal indvar222_601 : std_logic_vector(63 downto 0);
    signal indvar228_270 : std_logic_vector(63 downto 0);
    signal indvar231_189 : std_logic_vector(63 downto 0);
    signal indvar236_73 : std_logic_vector(63 downto 0);
    signal indvar_792 : std_logic_vector(63 downto 0);
    signal indvarx_xnext223_758 : std_logic_vector(63 downto 0);
    signal indvarx_xnext229_305 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_949 : std_logic_vector(63 downto 0);
    signal mul55_442 : std_logic_vector(63 downto 0);
    signal mul62_527 : std_logic_vector(63 downto 0);
    signal mul65_532 : std_logic_vector(63 downto 0);
    signal mul68_537 : std_logic_vector(63 downto 0);
    signal mul_437 : std_logic_vector(63 downto 0);
    signal ptr_deref_105_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_105_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_105_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_105_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_105_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_105_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_122_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_122_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_122_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_122_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_122_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_171_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_171_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_171_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_171_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_171_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_171_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_222_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_222_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_222_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_222_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_222_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_222_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_239_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_239_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_239_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_239_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_239_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_290_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_290_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_290_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_290_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_290_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_290_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_343_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_343_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_343_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_343_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_343_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_343_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_362_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_362_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_362_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_362_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_362_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_362_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_381_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_381_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_381_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_381_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_381_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_381_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_394_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_394_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_394_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_394_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_394_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_410_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_410_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_410_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_410_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_410_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_426_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_426_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_426_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_426_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_426_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_468_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_468_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_468_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_468_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_468_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_47_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_47_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_47_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_47_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_47_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_47_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_484_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_484_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_484_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_484_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_484_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_500_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_500_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_500_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_500_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_500_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_516_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_516_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_516_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_516_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_516_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_750_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_750_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_750_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_750_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_750_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_750_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_941_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_941_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_941_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_941_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_941_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_941_word_offset_0 : std_logic_vector(10 downto 0);
    signal sext192_542 : std_logic_vector(63 downto 0);
    signal sext_447 : std_logic_vector(63 downto 0);
    signal shl103_700 : std_logic_vector(63 downto 0);
    signal shl109_718 : std_logic_vector(63 downto 0);
    signal shl115_736 : std_logic_vector(63 downto 0);
    signal shl141_819 : std_logic_vector(63 downto 0);
    signal shl147_837 : std_logic_vector(63 downto 0);
    signal shl153_855 : std_logic_vector(63 downto 0);
    signal shl159_873 : std_logic_vector(63 downto 0);
    signal shl165_891 : std_logic_vector(63 downto 0);
    signal shl171_909 : std_logic_vector(63 downto 0);
    signal shl177_927 : std_logic_vector(63 downto 0);
    signal shl85_646 : std_logic_vector(63 downto 0);
    signal shl91_664 : std_logic_vector(63 downto 0);
    signal shl97_682 : std_logic_vector(63 downto 0);
    signal shl_628 : std_logic_vector(63 downto 0);
    signal shr132_776 : std_logic_vector(63 downto 0);
    signal shr_585 : std_logic_vector(63 downto 0);
    signal tmp12_240 : std_logic_vector(15 downto 0);
    signal tmp1_123 : std_logic_vector(15 downto 0);
    signal tmp233_230 : std_logic_vector(63 downto 0);
    signal tmp238_113 : std_logic_vector(63 downto 0);
    signal tmp2_92 : std_logic_vector(63 downto 0);
    signal tmp49_395 : std_logic_vector(15 downto 0);
    signal tmp4_202 : std_logic_vector(63 downto 0);
    signal tmp51_411 : std_logic_vector(15 downto 0);
    signal tmp53_427 : std_logic_vector(15 downto 0);
    signal tmp58_469 : std_logic_vector(15 downto 0);
    signal tmp60_485 : std_logic_vector(15 downto 0);
    signal tmp63_501 : std_logic_vector(15 downto 0);
    signal tmp66_517 : std_logic_vector(15 downto 0);
    signal tmp6_782 : std_logic_vector(0 downto 0);
    signal tmp_591 : std_logic_vector(0 downto 0);
    signal type_cast_111_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_131_wire : std_logic_vector(31 downto 0);
    signal type_cast_133_wire : std_logic_vector(31 downto 0);
    signal type_cast_153_wire : std_logic_vector(15 downto 0);
    signal type_cast_160_wire : std_logic_vector(15 downto 0);
    signal type_cast_162_wire : std_logic_vector(15 downto 0);
    signal type_cast_177_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_192_wire : std_logic_vector(63 downto 0);
    signal type_cast_195_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_200_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_228_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_247_wire : std_logic_vector(31 downto 0);
    signal type_cast_249_wire : std_logic_vector(31 downto 0);
    signal type_cast_274_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_276_wire : std_logic_vector(63 downto 0);
    signal type_cast_280_wire : std_logic_vector(15 downto 0);
    signal type_cast_282_wire : std_logic_vector(15 downto 0);
    signal type_cast_303_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_309_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_322_wire : std_logic_vector(15 downto 0);
    signal type_cast_435_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_451_wire : std_logic_vector(63 downto 0);
    signal type_cast_454_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_525_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_53_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_545_wire : std_logic_vector(63 downto 0);
    signal type_cast_548_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_555_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_570_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_583_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_589_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_596_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_605_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_607_wire : std_logic_vector(63 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_644_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_662_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_680_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_698_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_716_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_734_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_76_wire : std_logic_vector(63 downto 0);
    signal type_cast_774_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_780_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_787_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_798_wire : std_logic_vector(63 downto 0);
    signal type_cast_79_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_817_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_835_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_83_wire : std_logic_vector(15 downto 0);
    signal type_cast_853_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_85_wire : std_logic_vector(15 downto 0);
    signal type_cast_871_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_889_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_907_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_90_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_925_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_947_wire_constant : std_logic_vector(63 downto 0);
    signal umax7_789 : std_logic_vector(63 downto 0);
    signal umax_598 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_padding_324_word_address_0 <= "0";
    array_obj_ref_101_constant_part_of_offset <= "0000011";
    array_obj_ref_101_offset_scale_factor_0 <= "1000000";
    array_obj_ref_101_offset_scale_factor_1 <= "0000001";
    array_obj_ref_101_resized_base_address <= "0000000";
    array_obj_ref_211_constant_part_of_offset <= "0000011";
    array_obj_ref_211_offset_scale_factor_0 <= "1000000";
    array_obj_ref_211_offset_scale_factor_1 <= "0000001";
    array_obj_ref_211_resized_base_address <= "0000000";
    array_obj_ref_286_offset_scale_factor_0 <= "1";
    array_obj_ref_286_resized_base_address <= "0";
    array_obj_ref_613_constant_part_of_offset <= "00000000000000";
    array_obj_ref_613_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_613_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_613_resized_base_address <= "00000000000000";
    array_obj_ref_804_constant_part_of_offset <= "00000010001";
    array_obj_ref_804_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_804_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_804_resized_base_address <= "00000000000";
    iNsTr_13_119 <= "00000000000000000000000000000010";
    iNsTr_1_45 <= "00000000000000000000000000000010";
    iNsTr_21_236 <= "00000000000000000000000000000010";
    iNsTr_26_341 <= "00000000000000000000000000000011";
    iNsTr_29_360 <= "00000000000000000000000000000100";
    iNsTr_32_379 <= "00000000000000000000000000000101";
    iNsTr_34_391 <= "00000000000000000000000000000011";
    iNsTr_35_407 <= "00000000000000000000000000000100";
    iNsTr_36_423 <= "00000000000000000000000000000101";
    iNsTr_37_465 <= "00000000000000000000000000000011";
    iNsTr_38_481 <= "00000000000000000000000000000100";
    iNsTr_39_497 <= "00000000000000000000000000000101";
    iNsTr_40_513 <= "00000000000000000000000000000110";
    iNsTr_5_169 <= "00000000000000000000000000000010";
    ptr_deref_105_word_offset_0 <= "0000000";
    ptr_deref_122_word_offset_0 <= "0000000";
    ptr_deref_171_word_offset_0 <= "0000000";
    ptr_deref_222_word_offset_0 <= "0000000";
    ptr_deref_239_word_offset_0 <= "0000000";
    ptr_deref_290_word_offset_0 <= "0";
    ptr_deref_343_word_offset_0 <= "0000000";
    ptr_deref_362_word_offset_0 <= "0000000";
    ptr_deref_381_word_offset_0 <= "0000000";
    ptr_deref_394_word_offset_0 <= "0000000";
    ptr_deref_410_word_offset_0 <= "0000000";
    ptr_deref_426_word_offset_0 <= "0000000";
    ptr_deref_468_word_offset_0 <= "0000000";
    ptr_deref_47_word_offset_0 <= "0000000";
    ptr_deref_484_word_offset_0 <= "0000000";
    ptr_deref_500_word_offset_0 <= "0000000";
    ptr_deref_516_word_offset_0 <= "0000000";
    ptr_deref_750_word_offset_0 <= "00000000000000";
    ptr_deref_941_word_offset_0 <= "00000000000";
    type_cast_111_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_177_wire_constant <= "0000000000000000";
    type_cast_195_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_200_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_228_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_274_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_303_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_309_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_435_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_454_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_525_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_53_wire_constant <= "00000000";
    type_cast_548_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_555_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_570_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_583_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_589_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_596_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_605_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_626_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_644_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_662_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_680_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_698_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_716_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_734_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_756_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_774_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_780_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_787_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_796_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_79_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_817_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_835_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_853_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_871_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_889_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_907_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_90_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_925_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_947_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_150: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_153_wire;
      req(0) <= phi_stmt_150_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_150",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_150_ack_0,
          idata => idata,
          odata => conv5x_xlcssa1_150,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_150
    phi_stmt_157: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_160_wire & type_cast_162_wire;
      req <= phi_stmt_157_req_0 & phi_stmt_157_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_157",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_157_ack_0,
          idata => idata,
          odata => conv5x_xlcssa_157,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_157
    phi_stmt_189: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_192_wire & type_cast_195_wire_constant;
      req <= phi_stmt_189_req_0 & phi_stmt_189_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_189",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_189_ack_0,
          idata => idata,
          odata => indvar231_189,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_189
    phi_stmt_270: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_274_wire_constant & type_cast_276_wire;
      req <= phi_stmt_270_req_0 & phi_stmt_270_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_270",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_270_ack_0,
          idata => idata,
          odata => indvar228_270,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_270
    phi_stmt_277: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_280_wire & type_cast_282_wire;
      req <= phi_stmt_277_req_0 & phi_stmt_277_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_277",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_277_ack_0,
          idata => idata,
          odata => conv32206_277,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_277
    phi_stmt_319: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_322_wire;
      req(0) <= phi_stmt_319_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_319",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_319_ack_0,
          idata => idata,
          odata => conv32x_xlcssa_319,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_319
    phi_stmt_601: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_605_wire_constant & type_cast_607_wire;
      req <= phi_stmt_601_req_0 & phi_stmt_601_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_601",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_601_ack_0,
          idata => idata,
          odata => indvar222_601,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_601
    phi_stmt_73: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_76_wire & type_cast_79_wire_constant;
      req <= phi_stmt_73_req_0 & phi_stmt_73_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_73",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_73_ack_0,
          idata => idata,
          odata => indvar236_73,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_73
    phi_stmt_792: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_796_wire_constant & type_cast_798_wire;
      req <= phi_stmt_792_req_0 & phi_stmt_792_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_792",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_792_ack_0,
          idata => idata,
          odata => indvar_792,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_792
    phi_stmt_80: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_83_wire & type_cast_85_wire;
      req <= phi_stmt_80_req_0 & phi_stmt_80_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_80",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_80_ack_0,
          idata => idata,
          odata => conv5219_80,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_80
    -- flow-through select operator MUX_597_inst
    umax_598 <= shr_585 when (tmp_591(0) /=  '0') else type_cast_596_wire_constant;
    -- flow-through select operator MUX_788_inst
    umax7_789 <= shr132_776 when (tmp6_782(0) /=  '0') else type_cast_787_wire_constant;
    addr_of_102_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_102_final_reg_req_0;
      addr_of_102_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_102_final_reg_req_1;
      addr_of_102_final_reg_ack_1<= rack(0);
      addr_of_102_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_102_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_101_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_212_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_212_final_reg_req_0;
      addr_of_212_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_212_final_reg_req_1;
      addr_of_212_final_reg_ack_1<= rack(0);
      addr_of_212_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_212_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_211_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx21_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_287_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_287_final_reg_req_0;
      addr_of_287_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_287_final_reg_req_1;
      addr_of_287_final_reg_ack_1<= rack(0);
      addr_of_287_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_287_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_286_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx35_288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_614_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_614_final_reg_req_0;
      addr_of_614_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_614_final_reg_req_1;
      addr_of_614_final_reg_ack_1<= rack(0);
      addr_of_614_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_614_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_613_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx123_615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_805_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_805_final_reg_req_0;
      addr_of_805_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_805_final_reg_req_1;
      addr_of_805_final_reg_ack_1<= rack(0);
      addr_of_805_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_805_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_804_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx185_806,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp1_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_131_inst
    process(inc_96) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := inc_96(31 downto 0);
      type_cast_131_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_133_inst
    process(conv2_127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv2_127(31 downto 0);
      type_cast_133_wire <= tmp_var; -- 
    end process;
    type_cast_141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_141_inst_req_0;
      type_cast_141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_141_inst_req_1;
      type_cast_141_inst_ack_1<= rack(0);
      type_cast_141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5_142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_153_inst_req_0;
      type_cast_153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_153_inst_req_1;
      type_cast_153_inst_ack_1<= rack(0);
      type_cast_153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_153_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_160_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_160_inst_req_0;
      type_cast_160_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_160_inst_req_1;
      type_cast_160_inst_ack_1<= rack(0);
      type_cast_160_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_160_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5217_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_160_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_162_inst_req_0;
      type_cast_162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_162_inst_req_1;
      type_cast_162_inst_ack_1<= rack(0);
      type_cast_162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5x_xlcssa1_150,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_162_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_192_inst_req_0;
      type_cast_192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_192_inst_req_1;
      type_cast_192_inst_ack_1<= rack(0);
      type_cast_192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp233_230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_192_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_205_inst_req_0;
      type_cast_205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_205_inst_req_1;
      type_cast_205_inst_ack_1<= rack(0);
      type_cast_205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_202,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc24_206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_219_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_219_inst_req_0;
      type_cast_219_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_219_inst_req_1;
      type_cast_219_inst_ack_1<= rack(0);
      type_cast_219_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_219_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call17_216,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_220,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_243_inst_req_0;
      type_cast_243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_243_inst_req_1;
      type_cast_243_inst_ack_1<= rack(0);
      type_cast_243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_240,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_247_inst
    process(inc24_206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := inc24_206(31 downto 0);
      type_cast_247_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_249_inst
    process(conv13_244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv13_244(31 downto 0);
      type_cast_249_wire <= tmp_var; -- 
    end process;
    type_cast_266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_266_inst_req_0;
      type_cast_266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_266_inst_req_1;
      type_cast_266_inst_ack_1<= rack(0);
      type_cast_266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31203_263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32204_267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_276_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_276_inst_req_0;
      type_cast_276_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_276_inst_req_1;
      type_cast_276_inst_ack_1<= rack(0);
      type_cast_276_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_276_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext229_305,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_276_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_280_inst_req_0;
      type_cast_280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_280_inst_req_1;
      type_cast_280_inst_ack_1<= rack(0);
      type_cast_280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv32204_267,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_280_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_282_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_282_inst_req_0;
      type_cast_282_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_282_inst_req_1;
      type_cast_282_inst_ack_1<= rack(0);
      type_cast_282_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_282_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv32_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_282_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_298_inst_req_0;
      type_cast_298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_298_inst_req_1;
      type_cast_298_inst_ack_1<= rack(0);
      type_cast_298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_295,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_322_inst_req_0;
      type_cast_322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_322_inst_req_1;
      type_cast_322_inst_ack_1<= rack(0);
      type_cast_322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv32_299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_322_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_332_inst_req_0;
      type_cast_332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_332_inst_req_1;
      type_cast_332_inst_ack_1<= rack(0);
      type_cast_332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_329,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_333,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_351_inst_req_0;
      type_cast_351_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_351_inst_req_1;
      type_cast_351_inst_ack_1<= rack(0);
      type_cast_351_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_351_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_348,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_352,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_370_inst_req_0;
      type_cast_370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_370_inst_req_1;
      type_cast_370_inst_ack_1<= rack(0);
      type_cast_370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_398_inst_req_0;
      type_cast_398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_398_inst_req_1;
      type_cast_398_inst_ack_1<= rack(0);
      type_cast_398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp49_395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_414_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_414_inst_req_0;
      type_cast_414_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_414_inst_req_1;
      type_cast_414_inst_ack_1<= rack(0);
      type_cast_414_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_414_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp51_411,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_415,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_430_inst_req_0;
      type_cast_430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_430_inst_req_1;
      type_cast_430_inst_ack_1<= rack(0);
      type_cast_430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp53_427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv54_431,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_451_inst
    process(sext_447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_447(63 downto 0);
      type_cast_451_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_456_inst
    process(ASHR_i64_i64_455_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_455_wire(63 downto 0);
      conv56_457 <= tmp_var; -- 
    end process;
    type_cast_472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_472_inst_req_0;
      type_cast_472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_472_inst_req_1;
      type_cast_472_inst_ack_1<= rack(0);
      type_cast_472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp58_469,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_488_inst_req_0;
      type_cast_488_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_488_inst_req_1;
      type_cast_488_inst_ack_1<= rack(0);
      type_cast_488_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp60_485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_504_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_504_inst_req_0;
      type_cast_504_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_504_inst_req_1;
      type_cast_504_inst_ack_1<= rack(0);
      type_cast_504_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_504_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp63_501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_505,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_520_inst_req_0;
      type_cast_520_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_520_inst_req_1;
      type_cast_520_inst_ack_1<= rack(0);
      type_cast_520_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_520_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp66_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_545_inst
    process(sext192_542) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext192_542(63 downto 0);
      type_cast_545_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_550_inst
    process(ASHR_i64_i64_549_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_549_wire(63 downto 0);
      conv69_551 <= tmp_var; -- 
    end process;
    type_cast_607_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_607_inst_req_0;
      type_cast_607_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_607_inst_req_1;
      type_cast_607_inst_ack_1<= rack(0);
      type_cast_607_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_607_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext223_758,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_607_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_621_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_621_inst_req_0;
      type_cast_621_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_621_inst_req_1;
      type_cast_621_inst_ack_1<= rack(0);
      type_cast_621_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_621_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call78_618,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_622,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_62_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_62_inst_req_0;
      type_cast_62_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_62_inst_req_1;
      type_cast_62_inst_ack_1<= rack(0);
      type_cast_62_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_62_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4216_59,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5217_63,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_634_inst_req_0;
      type_cast_634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_634_inst_req_1;
      type_cast_634_inst_ack_1<= rack(0);
      type_cast_634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call81_631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_635,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_652_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_652_inst_req_0;
      type_cast_652_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_652_inst_req_1;
      type_cast_652_inst_ack_1<= rack(0);
      type_cast_652_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_652_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call86_649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_653,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_670_inst_req_0;
      type_cast_670_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_670_inst_req_1;
      type_cast_670_inst_ack_1<= rack(0);
      type_cast_670_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_670_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_667,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_688_inst_req_0;
      type_cast_688_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_688_inst_req_1;
      type_cast_688_inst_ack_1<= rack(0);
      type_cast_688_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_688_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call98_685,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_689,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_706_inst_req_0;
      type_cast_706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_706_inst_req_1;
      type_cast_706_inst_ack_1<= rack(0);
      type_cast_706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call104_703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv106_707,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_724_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_724_inst_req_0;
      type_cast_724_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_724_inst_req_1;
      type_cast_724_inst_ack_1<= rack(0);
      type_cast_724_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_724_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_725,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_742_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_742_inst_req_0;
      type_cast_742_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_742_inst_req_1;
      type_cast_742_inst_ack_1<= rack(0);
      type_cast_742_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_742_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call116_739,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_743,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp238_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_76_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_798_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_798_inst_req_0;
      type_cast_798_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_798_inst_req_1;
      type_cast_798_inst_ack_1<= rack(0);
      type_cast_798_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_798_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_949,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_798_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_812_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_812_inst_req_0;
      type_cast_812_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_812_inst_req_1;
      type_cast_812_inst_ack_1<= rack(0);
      type_cast_812_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_812_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call138_809,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv139_813,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_825_inst_req_0;
      type_cast_825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_825_inst_req_1;
      type_cast_825_inst_ack_1<= rack(0);
      type_cast_825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call142_822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_83_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_83_inst_req_0;
      type_cast_83_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_83_inst_req_1;
      type_cast_83_inst_ack_1<= rack(0);
      type_cast_83_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_83_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5_142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_83_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_843_inst_req_0;
      type_cast_843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_843_inst_req_1;
      type_cast_843_inst_ack_1<= rack(0);
      type_cast_843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call148_840,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv150_844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_85_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_85_inst_req_0;
      type_cast_85_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_85_inst_req_1;
      type_cast_85_inst_ack_1<= rack(0);
      type_cast_85_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_85_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv5217_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_85_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_861_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_861_inst_req_0;
      type_cast_861_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_861_inst_req_1;
      type_cast_861_inst_ack_1<= rack(0);
      type_cast_861_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_861_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call154_858,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv156_862,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_879_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_879_inst_req_0;
      type_cast_879_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_879_inst_req_1;
      type_cast_879_inst_ack_1<= rack(0);
      type_cast_879_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_879_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call160_876,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv162_880,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_897_inst_req_0;
      type_cast_897_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_897_inst_req_1;
      type_cast_897_inst_ack_1<= rack(0);
      type_cast_897_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_897_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call166_894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv168_898,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_915_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_915_inst_req_0;
      type_cast_915_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_915_inst_req_1;
      type_cast_915_inst_ack_1<= rack(0);
      type_cast_915_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_915_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call172_912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv174_916,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_933_inst_req_0;
      type_cast_933_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_933_inst_req_1;
      type_cast_933_inst_ack_1<= rack(0);
      type_cast_933_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call178_930,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv180_934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp2_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_966_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_966_inst_req_0;
      type_cast_966_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_966_inst_req_1;
      type_cast_966_inst_ack_1<= rack(0);
      type_cast_966_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_966_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv56_457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_padding_324_gather_scatter
    process(conv32x_xlcssa_319) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv32x_xlcssa_319;
      ov(15 downto 0) := iv;
      STORE_padding_324_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_rename
    process(R_indvar236_100_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar236_100_resized;
      ov(6 downto 0) := iv;
      R_indvar236_100_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_resize
    process(indvar236_73) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar236_73;
      ov := iv(6 downto 0);
      R_indvar236_100_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_root_address_inst
    process(array_obj_ref_101_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_101_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_101_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_211_index_1_rename
    process(R_indvar231_210_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar231_210_resized;
      ov(6 downto 0) := iv;
      R_indvar231_210_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_211_index_1_resize
    process(indvar231_189) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar231_189;
      ov := iv(6 downto 0);
      R_indvar231_210_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_211_root_address_inst
    process(array_obj_ref_211_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_211_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_211_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_286_index_0_rename
    process(R_indvar228_285_resized) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar228_285_resized;
      ov(0 downto 0) := iv;
      R_indvar228_285_scaled <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_286_index_0_resize
    process(indvar228_270) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar228_270;
      ov := iv(0 downto 0);
      R_indvar228_285_resized <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_286_index_offset
    process(R_indvar228_285_scaled) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar228_285_scaled;
      ov(0 downto 0) := iv;
      array_obj_ref_286_final_offset <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_286_root_address_inst
    process(array_obj_ref_286_final_offset) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_286_final_offset;
      ov(0 downto 0) := iv;
      array_obj_ref_286_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_613_index_1_rename
    process(R_indvar222_612_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar222_612_resized;
      ov(13 downto 0) := iv;
      R_indvar222_612_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_613_index_1_resize
    process(indvar222_601) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar222_601;
      ov := iv(13 downto 0);
      R_indvar222_612_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_613_root_address_inst
    process(array_obj_ref_613_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_613_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_613_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_804_index_1_rename
    process(R_indvar_803_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_803_resized;
      ov(10 downto 0) := iv;
      R_indvar_803_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_804_index_1_resize
    process(indvar_792) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_792;
      ov := iv(10 downto 0);
      R_indvar_803_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_804_root_address_inst
    process(array_obj_ref_804_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_804_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_804_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_addr_0
    process(ptr_deref_105_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_105_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_105_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_base_resize
    process(arrayidx_103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_103;
      ov := iv(6 downto 0);
      ptr_deref_105_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_gather_scatter
    process(conv5219_80) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv5219_80;
      ov(15 downto 0) := iv;
      ptr_deref_105_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_root_address_inst
    process(ptr_deref_105_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_105_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_105_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_addr_0
    process(ptr_deref_122_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_122_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_base_resize
    process(iNsTr_13_119) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_13_119;
      ov := iv(6 downto 0);
      ptr_deref_122_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_gather_scatter
    process(ptr_deref_122_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_data_0;
      ov(15 downto 0) := iv;
      tmp1_123 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_root_address_inst
    process(ptr_deref_122_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_122_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_171_addr_0
    process(ptr_deref_171_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_171_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_171_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_171_base_resize
    process(iNsTr_5_169) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_169;
      ov := iv(6 downto 0);
      ptr_deref_171_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_171_gather_scatter
    process(conv5x_xlcssa_157) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv5x_xlcssa_157;
      ov(15 downto 0) := iv;
      ptr_deref_171_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_171_root_address_inst
    process(ptr_deref_171_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_171_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_171_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_222_addr_0
    process(ptr_deref_222_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_222_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_222_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_222_base_resize
    process(arrayidx21_213) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx21_213;
      ov := iv(6 downto 0);
      ptr_deref_222_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_222_gather_scatter
    process(conv18_220) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv18_220;
      ov(15 downto 0) := iv;
      ptr_deref_222_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_222_root_address_inst
    process(ptr_deref_222_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_222_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_222_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_239_addr_0
    process(ptr_deref_239_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_239_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_239_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_239_base_resize
    process(iNsTr_21_236) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_236;
      ov := iv(6 downto 0);
      ptr_deref_239_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_239_gather_scatter
    process(ptr_deref_239_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_239_data_0;
      ov(15 downto 0) := iv;
      tmp12_240 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_239_root_address_inst
    process(ptr_deref_239_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_239_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_239_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_290_addr_0
    process(ptr_deref_290_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_290_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_290_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_290_base_resize
    process(arrayidx35_288) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx35_288;
      ov := iv(0 downto 0);
      ptr_deref_290_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_290_gather_scatter
    process(conv32206_277) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv32206_277;
      ov(15 downto 0) := iv;
      ptr_deref_290_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_290_root_address_inst
    process(ptr_deref_290_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_290_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_290_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_addr_0
    process(ptr_deref_343_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_343_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_base_resize
    process(iNsTr_26_341) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_341;
      ov := iv(6 downto 0);
      ptr_deref_343_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_gather_scatter
    process(conv43_333) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv43_333;
      ov(15 downto 0) := iv;
      ptr_deref_343_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_root_address_inst
    process(ptr_deref_343_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_343_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_362_addr_0
    process(ptr_deref_362_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_362_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_362_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_362_base_resize
    process(iNsTr_29_360) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_29_360;
      ov := iv(6 downto 0);
      ptr_deref_362_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_362_gather_scatter
    process(conv45_352) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv45_352;
      ov(15 downto 0) := iv;
      ptr_deref_362_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_362_root_address_inst
    process(ptr_deref_362_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_362_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_362_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_addr_0
    process(ptr_deref_381_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_381_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_base_resize
    process(iNsTr_32_379) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_32_379;
      ov := iv(6 downto 0);
      ptr_deref_381_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_gather_scatter
    process(conv47_371) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv47_371;
      ov(15 downto 0) := iv;
      ptr_deref_381_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_root_address_inst
    process(ptr_deref_381_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_381_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_addr_0
    process(ptr_deref_394_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_394_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_base_resize
    process(iNsTr_34_391) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_391;
      ov := iv(6 downto 0);
      ptr_deref_394_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_gather_scatter
    process(ptr_deref_394_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_data_0;
      ov(15 downto 0) := iv;
      tmp49_395 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_394_root_address_inst
    process(ptr_deref_394_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_394_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_394_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_410_addr_0
    process(ptr_deref_410_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_410_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_410_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_410_base_resize
    process(iNsTr_35_407) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_35_407;
      ov := iv(6 downto 0);
      ptr_deref_410_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_410_gather_scatter
    process(ptr_deref_410_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_410_data_0;
      ov(15 downto 0) := iv;
      tmp51_411 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_410_root_address_inst
    process(ptr_deref_410_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_410_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_410_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_addr_0
    process(ptr_deref_426_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_426_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_base_resize
    process(iNsTr_36_423) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_36_423;
      ov := iv(6 downto 0);
      ptr_deref_426_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_gather_scatter
    process(ptr_deref_426_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_data_0;
      ov(15 downto 0) := iv;
      tmp53_427 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_426_root_address_inst
    process(ptr_deref_426_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_426_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_426_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_addr_0
    process(ptr_deref_468_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_468_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_base_resize
    process(iNsTr_37_465) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_465;
      ov := iv(6 downto 0);
      ptr_deref_468_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_gather_scatter
    process(ptr_deref_468_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_data_0;
      ov(15 downto 0) := iv;
      tmp58_469 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_468_root_address_inst
    process(ptr_deref_468_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_468_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_468_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_addr_0
    process(ptr_deref_47_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_47_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_47_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_base_resize
    process(iNsTr_1_45) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_45;
      ov := iv(6 downto 0);
      ptr_deref_47_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_gather_scatter
    process(conv_39) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_39;
      ov(15 downto 0) := iv;
      ptr_deref_47_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_root_address_inst
    process(ptr_deref_47_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_47_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_47_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_484_addr_0
    process(ptr_deref_484_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_484_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_484_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_484_base_resize
    process(iNsTr_38_481) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_481;
      ov := iv(6 downto 0);
      ptr_deref_484_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_484_gather_scatter
    process(ptr_deref_484_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_484_data_0;
      ov(15 downto 0) := iv;
      tmp60_485 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_484_root_address_inst
    process(ptr_deref_484_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_484_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_484_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_addr_0
    process(ptr_deref_500_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_500_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_500_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_base_resize
    process(iNsTr_39_497) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_39_497;
      ov := iv(6 downto 0);
      ptr_deref_500_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_gather_scatter
    process(ptr_deref_500_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_500_data_0;
      ov(15 downto 0) := iv;
      tmp63_501 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_500_root_address_inst
    process(ptr_deref_500_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_500_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_500_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_516_addr_0
    process(ptr_deref_516_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_516_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_516_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_516_base_resize
    process(iNsTr_40_513) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_513;
      ov := iv(6 downto 0);
      ptr_deref_516_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_516_gather_scatter
    process(ptr_deref_516_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_516_data_0;
      ov(15 downto 0) := iv;
      tmp66_517 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_516_root_address_inst
    process(ptr_deref_516_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_516_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_516_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_750_addr_0
    process(ptr_deref_750_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_750_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_750_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_750_base_resize
    process(arrayidx123_615) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx123_615;
      ov := iv(13 downto 0);
      ptr_deref_750_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_750_gather_scatter
    process(add119_748) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add119_748;
      ov(63 downto 0) := iv;
      ptr_deref_750_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_750_root_address_inst
    process(ptr_deref_750_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_750_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_750_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_addr_0
    process(ptr_deref_941_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_941_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_941_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_base_resize
    process(arrayidx185_806) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx185_806;
      ov := iv(10 downto 0);
      ptr_deref_941_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_gather_scatter
    process(add181_939) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add181_939;
      ov(63 downto 0) := iv;
      ptr_deref_941_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_root_address_inst
    process(ptr_deref_941_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_941_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_941_root_address <= ov(10 downto 0);
      --
    end process;
    if_stmt_143_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_135;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_143_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_143_branch_req_0,
          ack0 => if_stmt_143_branch_ack_0,
          ack1 => if_stmt_143_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_180_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp14210_179;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_180_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_180_branch_req_0,
          ack0 => if_stmt_180_branch_ack_0,
          ack1 => if_stmt_180_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_252_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp14_251;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_252_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_252_branch_req_0,
          ack0 => if_stmt_252_branch_ack_0,
          ack1 => if_stmt_252_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_312_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond9_311;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_312_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_312_branch_req_0,
          ack0 => if_stmt_312_branch_ack_0,
          ack1 => if_stmt_312_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_558_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp74199_557;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_558_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_558_branch_req_0,
          ack0 => if_stmt_558_branch_ack_0,
          ack1 => if_stmt_558_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_573_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp133195_572;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_573_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_573_branch_req_0,
          ack0 => if_stmt_573_branch_ack_0,
          ack1 => if_stmt_573_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_64_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp215_56;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_64_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_64_branch_req_0,
          ack0 => if_stmt_64_branch_ack_0,
          ack1 => if_stmt_64_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_764_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_763;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_764_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_764_branch_req_0,
          ack0 => if_stmt_764_branch_ack_0,
          ack1 => if_stmt_764_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_955_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond8_954;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_955_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_955_branch_req_0,
          ack0 => if_stmt_955_branch_ack_0,
          ack1 => if_stmt_955_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_112_inst
    process(indvar236_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar236_73, type_cast_111_wire_constant, tmp_var);
      tmp238_113 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_201_inst
    process(indvar231_189) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar231_189, type_cast_200_wire_constant, tmp_var);
      tmp4_202 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_229_inst
    process(indvar231_189) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar231_189, type_cast_228_wire_constant, tmp_var);
      tmp233_230 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_304_inst
    process(indvar228_270) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar228_270, type_cast_303_wire_constant, tmp_var);
      indvarx_xnext229_305 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_757_inst
    process(indvar222_601) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar222_601, type_cast_756_wire_constant, tmp_var);
      indvarx_xnext223_758 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_91_inst
    process(indvar236_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar236_73, type_cast_90_wire_constant, tmp_var);
      tmp2_92 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_948_inst
    process(indvar_792) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_792, type_cast_947_wire_constant, tmp_var);
      indvarx_xnext_949 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_455_inst
    process(type_cast_451_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_451_wire, type_cast_454_wire_constant, tmp_var);
      ASHR_i64_i64_455_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_549_inst
    process(type_cast_545_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_545_wire, type_cast_548_wire_constant, tmp_var);
      ASHR_i64_i64_549_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_178_inst
    process(conv5x_xlcssa_157) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv5x_xlcssa_157, type_cast_177_wire_constant, tmp_var);
      cmp14210_179 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_310_inst
    process(indvarx_xnext229_305) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext229_305, type_cast_309_wire_constant, tmp_var);
      exitcond9_311 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_762_inst
    process(indvarx_xnext223_758, umax_598) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext223_758, umax_598, tmp_var);
      exitcond_763 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_953_inst
    process(indvarx_xnext_949, umax7_789) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_949, umax7_789, tmp_var);
      exitcond8_954 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_54_inst
    process(call_35) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(call_35, type_cast_53_wire_constant, tmp_var);
      cmp215_56 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_584_inst
    process(conv56_457) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv56_457, type_cast_583_wire_constant, tmp_var);
      shr_585 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_775_inst
    process(conv69_551) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv69_551, type_cast_774_wire_constant, tmp_var);
      shr132_776 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_441_inst
    process(mul_437, conv52_415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_437, conv52_415, tmp_var);
      mul55_442 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_446_inst
    process(mul55_442, conv54_431) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul55_442, conv54_431, tmp_var);
      sext_447 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_531_inst
    process(mul62_527, conv61_489) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul62_527, conv61_489, tmp_var);
      mul65_532 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_536_inst
    process(mul65_532, conv64_505) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul65_532, conv64_505, tmp_var);
      mul68_537 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_541_inst
    process(mul68_537, conv67_521) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul68_537, conv67_521, tmp_var);
      sext192_542 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_639_inst
    process(shl_628, conv83_635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_628, conv83_635, tmp_var);
      add_640 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_657_inst
    process(shl85_646, conv88_653) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl85_646, conv88_653, tmp_var);
      add89_658 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_675_inst
    process(shl91_664, conv94_671) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl91_664, conv94_671, tmp_var);
      add95_676 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_693_inst
    process(shl97_682, conv100_689) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl97_682, conv100_689, tmp_var);
      add101_694 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_711_inst
    process(shl103_700, conv106_707) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl103_700, conv106_707, tmp_var);
      add107_712 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_729_inst
    process(shl109_718, conv112_725) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl109_718, conv112_725, tmp_var);
      add113_730 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_747_inst
    process(shl115_736, conv118_743) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl115_736, conv118_743, tmp_var);
      add119_748 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_830_inst
    process(shl141_819, conv144_826) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl141_819, conv144_826, tmp_var);
      add145_831 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_848_inst
    process(shl147_837, conv150_844) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl147_837, conv150_844, tmp_var);
      add151_849 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_866_inst
    process(shl153_855, conv156_862) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl153_855, conv156_862, tmp_var);
      add157_867 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_884_inst
    process(shl159_873, conv162_880) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl159_873, conv162_880, tmp_var);
      add163_885 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_902_inst
    process(shl165_891, conv168_898) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl165_891, conv168_898, tmp_var);
      add169_903 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_920_inst
    process(shl171_909, conv174_916) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl171_909, conv174_916, tmp_var);
      add175_921 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_938_inst
    process(shl177_927, conv180_934) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl177_927, conv180_934, tmp_var);
      add181_939 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_436_inst
    process(conv50_399) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv50_399, type_cast_435_wire_constant, tmp_var);
      mul_437 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_526_inst
    process(conv59_473) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_473, type_cast_525_wire_constant, tmp_var);
      mul62_527 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_627_inst
    process(conv79_622) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv79_622, type_cast_626_wire_constant, tmp_var);
      shl_628 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_645_inst
    process(add_640) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_640, type_cast_644_wire_constant, tmp_var);
      shl85_646 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_663_inst
    process(add89_658) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add89_658, type_cast_662_wire_constant, tmp_var);
      shl91_664 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_681_inst
    process(add95_676) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add95_676, type_cast_680_wire_constant, tmp_var);
      shl97_682 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_699_inst
    process(add101_694) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add101_694, type_cast_698_wire_constant, tmp_var);
      shl103_700 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_717_inst
    process(add107_712) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add107_712, type_cast_716_wire_constant, tmp_var);
      shl109_718 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_735_inst
    process(add113_730) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add113_730, type_cast_734_wire_constant, tmp_var);
      shl115_736 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_818_inst
    process(conv139_813) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv139_813, type_cast_817_wire_constant, tmp_var);
      shl141_819 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_836_inst
    process(add145_831) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add145_831, type_cast_835_wire_constant, tmp_var);
      shl147_837 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_854_inst
    process(add151_849) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add151_849, type_cast_853_wire_constant, tmp_var);
      shl153_855 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_872_inst
    process(add157_867) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add157_867, type_cast_871_wire_constant, tmp_var);
      shl159_873 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_890_inst
    process(add163_885) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add163_885, type_cast_889_wire_constant, tmp_var);
      shl165_891 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_908_inst
    process(add169_903) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add169_903, type_cast_907_wire_constant, tmp_var);
      shl171_909 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_926_inst
    process(add175_921) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add175_921, type_cast_925_wire_constant, tmp_var);
      shl177_927 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_134_inst
    process(type_cast_131_wire, type_cast_133_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_131_wire, type_cast_133_wire, tmp_var);
      cmp_135 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_250_inst
    process(type_cast_247_wire, type_cast_249_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_247_wire, type_cast_249_wire, tmp_var);
      cmp14_251 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_556_inst
    process(conv56_457) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv56_457, type_cast_555_wire_constant, tmp_var);
      cmp74199_557 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_571_inst
    process(conv69_551) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv69_551, type_cast_570_wire_constant, tmp_var);
      cmp133195_572 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_590_inst
    process(shr_585) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_585, type_cast_589_wire_constant, tmp_var);
      tmp_591 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_781_inst
    process(shr132_776) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr132_776, type_cast_780_wire_constant, tmp_var);
      tmp6_782 <= tmp_var; --
    end process;
    -- shared split operator group (57) : array_obj_ref_101_index_offset 
    ApIntAdd_group_57: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar236_100_scaled;
      array_obj_ref_101_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_101_index_offset_req_0;
      array_obj_ref_101_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_101_index_offset_req_1;
      array_obj_ref_101_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_57_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_57_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_57",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000011",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : array_obj_ref_211_index_offset 
    ApIntAdd_group_58: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar231_210_scaled;
      array_obj_ref_211_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_211_index_offset_req_0;
      array_obj_ref_211_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_211_index_offset_req_1;
      array_obj_ref_211_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_58_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_58_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_58",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000011",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : array_obj_ref_613_index_offset 
    ApIntAdd_group_59: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar222_612_scaled;
      array_obj_ref_613_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_613_index_offset_req_0;
      array_obj_ref_613_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_613_index_offset_req_1;
      array_obj_ref_613_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_59_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_59_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_59",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : array_obj_ref_804_index_offset 
    ApIntAdd_group_60: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_803_scaled;
      array_obj_ref_804_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_804_index_offset_req_0;
      array_obj_ref_804_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_804_index_offset_req_1;
      array_obj_ref_804_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_60_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_60_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_60",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000010001",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared load operator group (0) : ptr_deref_122_load_0 ptr_deref_394_load_0 ptr_deref_410_load_0 ptr_deref_426_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_122_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_394_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_410_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_426_load_0_req_0;
      ptr_deref_122_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_394_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_410_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_426_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_122_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_394_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_410_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_426_load_0_req_1;
      ptr_deref_122_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_394_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_410_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_426_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_122_word_address_0 & ptr_deref_394_word_address_0 & ptr_deref_410_word_address_0 & ptr_deref_426_word_address_0;
      ptr_deref_122_data_0 <= data_out(63 downto 48);
      ptr_deref_394_data_0 <= data_out(47 downto 32);
      ptr_deref_410_data_0 <= data_out(31 downto 16);
      ptr_deref_426_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(15 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_239_load_0 ptr_deref_468_load_0 ptr_deref_484_load_0 ptr_deref_500_load_0 ptr_deref_516_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(34 downto 0);
      signal data_out: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= ptr_deref_239_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_468_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_484_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_500_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_516_load_0_req_0;
      ptr_deref_239_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_468_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_484_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_500_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_516_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= ptr_deref_239_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_468_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_484_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_500_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_516_load_0_req_1;
      ptr_deref_239_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_468_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_484_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_500_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_516_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_239_word_address_0 & ptr_deref_468_word_address_0 & ptr_deref_484_word_address_0 & ptr_deref_500_word_address_0 & ptr_deref_516_word_address_0;
      ptr_deref_239_data_0 <= data_out(79 downto 64);
      ptr_deref_468_data_0 <= data_out(63 downto 48);
      ptr_deref_484_data_0 <= data_out(47 downto 32);
      ptr_deref_500_data_0 <= data_out(31 downto 16);
      ptr_deref_516_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 16,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(15 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared store operator group (0) : STORE_padding_324_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_padding_324_store_0_req_0;
      STORE_padding_324_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_padding_324_store_0_req_1;
      STORE_padding_324_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_padding_324_word_address_0;
      data_in <= STORE_padding_324_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(15 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_47_store_0 ptr_deref_105_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_47_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_105_store_0_req_0;
      ptr_deref_47_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_105_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_47_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_105_store_0_req_1;
      ptr_deref_47_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_105_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_47_word_address_0 & ptr_deref_105_word_address_0;
      data_in <= ptr_deref_47_data_0 & ptr_deref_105_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(6 downto 0),
          mdata => memory_space_0_sr_data(15 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_222_store_0 ptr_deref_171_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_222_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_171_store_0_req_0;
      ptr_deref_222_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_171_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_222_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_171_store_0_req_1;
      ptr_deref_222_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_171_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_222_word_address_0 & ptr_deref_171_word_address_0;
      data_in <= ptr_deref_222_data_0 & ptr_deref_171_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(15 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_290_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_290_store_0_req_0;
      ptr_deref_290_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_290_store_0_req_1;
      ptr_deref_290_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_290_word_address_0;
      data_in <= ptr_deref_290_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_343_store_0 ptr_deref_362_store_0 ptr_deref_381_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_343_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_362_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_381_store_0_req_0;
      ptr_deref_343_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_362_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_381_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_343_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_362_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_381_store_0_req_1;
      ptr_deref_343_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_362_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_381_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup4_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_343_word_address_0 & ptr_deref_362_word_address_0 & ptr_deref_381_word_address_0;
      data_in <= ptr_deref_343_data_0 & ptr_deref_362_data_0 & ptr_deref_381_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 7,
        data_width => 16,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(15 downto 0),
          mtag => memory_space_2_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_750_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_750_store_0_req_0;
      ptr_deref_750_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_750_store_0_req_1;
      ptr_deref_750_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_750_word_address_0;
      data_in <= ptr_deref_750_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_941_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_941_store_0_req_0;
      ptr_deref_941_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_941_store_0_req_1;
      ptr_deref_941_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_941_word_address_0;
      data_in <= ptr_deref_941_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(10 downto 0),
          mdata => memory_space_4_sr_data(63 downto 0),
          mtag => memory_space_4_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_808_inst RPIPE_ConvTranspose_input_pipe_821_inst RPIPE_ConvTranspose_input_pipe_702_inst RPIPE_ConvTranspose_input_pipe_720_inst RPIPE_ConvTranspose_input_pipe_929_inst RPIPE_ConvTranspose_input_pipe_839_inst RPIPE_ConvTranspose_input_pipe_857_inst RPIPE_ConvTranspose_input_pipe_738_inst RPIPE_ConvTranspose_input_pipe_875_inst RPIPE_ConvTranspose_input_pipe_893_inst RPIPE_ConvTranspose_input_pipe_58_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_684_inst RPIPE_ConvTranspose_input_pipe_911_inst RPIPE_ConvTranspose_input_pipe_648_inst RPIPE_ConvTranspose_input_pipe_617_inst RPIPE_ConvTranspose_input_pipe_630_inst RPIPE_ConvTranspose_input_pipe_137_inst RPIPE_ConvTranspose_input_pipe_215_inst RPIPE_ConvTranspose_input_pipe_262_inst RPIPE_ConvTranspose_input_pipe_666_inst RPIPE_ConvTranspose_input_pipe_294_inst RPIPE_ConvTranspose_input_pipe_328_inst RPIPE_ConvTranspose_input_pipe_347_inst RPIPE_ConvTranspose_input_pipe_366_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(199 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 24 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 24 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 24 downto 0);
      signal guard_vector : std_logic_vector( 24 downto 0);
      constant outBUFs : IntegerArray(24 downto 0) := (24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(24 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false);
      constant guardBuffering: IntegerArray(24 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2);
      -- 
    begin -- 
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_808_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_821_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_702_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_720_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_929_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_839_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_857_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_738_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_875_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_893_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_58_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_684_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_911_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_648_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_617_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_630_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_137_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_215_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_262_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_666_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_294_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_328_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_347_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_808_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_821_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_702_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_720_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_929_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_839_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_857_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_738_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_875_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_893_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_58_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_684_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_911_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_648_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_617_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_630_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_137_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_215_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_262_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_666_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_294_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_328_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_347_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_808_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_821_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_702_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_720_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_929_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_839_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_857_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_738_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_875_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_893_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_58_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_684_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_911_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_648_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_617_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_630_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_137_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_215_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_262_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_666_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_294_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_328_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_347_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_808_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_821_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_702_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_720_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_929_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_839_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_857_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_738_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_875_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_893_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_58_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_684_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_911_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_648_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_617_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_630_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_137_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_215_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_262_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_666_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_294_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_328_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_347_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      call138_809 <= data_out(199 downto 192);
      call142_822 <= data_out(191 downto 184);
      call104_703 <= data_out(183 downto 176);
      call110_721 <= data_out(175 downto 168);
      call178_930 <= data_out(167 downto 160);
      call148_840 <= data_out(159 downto 152);
      call154_858 <= data_out(151 downto 144);
      call116_739 <= data_out(143 downto 136);
      call160_876 <= data_out(135 downto 128);
      call166_894 <= data_out(127 downto 120);
      call4216_59 <= data_out(119 downto 112);
      call_35 <= data_out(111 downto 104);
      call98_685 <= data_out(103 downto 96);
      call172_912 <= data_out(95 downto 88);
      call86_649 <= data_out(87 downto 80);
      call78_618 <= data_out(79 downto 72);
      call81_631 <= data_out(71 downto 64);
      call4_138 <= data_out(63 downto 56);
      call17_216 <= data_out(55 downto 48);
      call31203_263 <= data_out(47 downto 40);
      call92_667 <= data_out(39 downto 32);
      call31_295 <= data_out(31 downto 24);
      call42_329 <= data_out(23 downto 16);
      call44_348 <= data_out(15 downto 8);
      call46_367 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 25, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 25,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(99 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(3 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(3 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(55 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(75 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(3 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 21),
      memory_space_0_lr_tag => memory_space_0_lr_tag(83 downto 63),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 48),
      memory_space_0_lc_tag => memory_space_0_lc_tag(11 downto 9),
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 21),
      memory_space_1_lr_tag => memory_space_1_lr_tag(83 downto 63),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 48),
      memory_space_1_lc_tag => memory_space_1_lc_tag(11 downto 9),
      memory_space_2_lr_req => memory_space_2_lr_req(4 downto 4),
      memory_space_2_lr_ack => memory_space_2_lr_ack(4 downto 4),
      memory_space_2_lr_addr => memory_space_2_lr_addr(34 downto 28),
      memory_space_2_lr_tag => memory_space_2_lr_tag(99 downto 80),
      memory_space_2_lc_req => memory_space_2_lc_req(4 downto 4),
      memory_space_2_lc_ack => memory_space_2_lc_ack(4 downto 4),
      memory_space_2_lc_data => memory_space_2_lc_data(79 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(9 downto 8),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(55 downto 42),
      memory_space_3_lr_tag => memory_space_3_lr_tag(75 downto 57),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(255 downto 192),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 3),
      memory_space_6_lr_req => memory_space_6_lr_req(3 downto 3),
      memory_space_6_lr_ack => memory_space_6_lr_ack(3 downto 3),
      memory_space_6_lr_addr => memory_space_6_lr_addr(3 downto 3),
      memory_space_6_lr_tag => memory_space_6_lr_tag(75 downto 57),
      memory_space_6_lc_req => memory_space_6_lc_req(3 downto 3),
      memory_space_6_lc_ack => memory_space_6_lc_ack(3 downto 3),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 48),
      memory_space_6_lc_tag => memory_space_6_lc_tag(3 downto 3),
      memory_space_7_lr_req => memory_space_7_lr_req(3 downto 3),
      memory_space_7_lr_ack => memory_space_7_lr_ack(3 downto 3),
      memory_space_7_lr_addr => memory_space_7_lr_addr(3 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(79 downto 60),
      memory_space_7_lc_req => memory_space_7_lc_req(3 downto 3),
      memory_space_7_lc_ack => memory_space_7_lc_ack(3 downto 3),
      memory_space_7_lc_data => memory_space_7_lc_data(63 downto 48),
      memory_space_7_lc_tag => memory_space_7_lc_tag(7 downto 6),
      memory_space_5_sr_req => memory_space_5_sr_req(3 downto 3),
      memory_space_5_sr_ack => memory_space_5_sr_ack(3 downto 3),
      memory_space_5_sr_addr => memory_space_5_sr_addr(55 downto 42),
      memory_space_5_sr_data => memory_space_5_sr_data(255 downto 192),
      memory_space_5_sr_tag => memory_space_5_sr_tag(75 downto 57),
      memory_space_5_sc_req => memory_space_5_sc_req(3 downto 3),
      memory_space_5_sc_ack => memory_space_5_sc_ack(3 downto 3),
      memory_space_5_sc_tag => memory_space_5_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(20 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(62 downto 42),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(47 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(8 downto 6),
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(20 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(62 downto 42),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(47 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(8 downto 6),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(20 downto 14),
      memory_space_2_lr_tag => memory_space_2_lr_tag(59 downto 40),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(47 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 4),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(41 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(56 downto 38),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(191 downto 128),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 2),
      memory_space_6_lr_req => memory_space_6_lr_req(2 downto 2),
      memory_space_6_lr_ack => memory_space_6_lr_ack(2 downto 2),
      memory_space_6_lr_addr => memory_space_6_lr_addr(2 downto 2),
      memory_space_6_lr_tag => memory_space_6_lr_tag(56 downto 38),
      memory_space_6_lc_req => memory_space_6_lc_req(2 downto 2),
      memory_space_6_lc_ack => memory_space_6_lc_ack(2 downto 2),
      memory_space_6_lc_data => memory_space_6_lc_data(47 downto 32),
      memory_space_6_lc_tag => memory_space_6_lc_tag(2 downto 2),
      memory_space_7_lr_req => memory_space_7_lr_req(2 downto 2),
      memory_space_7_lr_ack => memory_space_7_lr_ack(2 downto 2),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 2),
      memory_space_7_lr_tag => memory_space_7_lr_tag(59 downto 40),
      memory_space_7_lc_req => memory_space_7_lc_req(2 downto 2),
      memory_space_7_lc_ack => memory_space_7_lc_ack(2 downto 2),
      memory_space_7_lc_data => memory_space_7_lc_data(47 downto 32),
      memory_space_7_lc_tag => memory_space_7_lc_tag(5 downto 4),
      memory_space_5_sr_req => memory_space_5_sr_req(2 downto 2),
      memory_space_5_sr_ack => memory_space_5_sr_ack(2 downto 2),
      memory_space_5_sr_addr => memory_space_5_sr_addr(41 downto 28),
      memory_space_5_sr_data => memory_space_5_sr_data(191 downto 128),
      memory_space_5_sr_tag => memory_space_5_sr_tag(56 downto 38),
      memory_space_5_sc_req => memory_space_5_sc_req(2 downto 2),
      memory_space_5_sc_ack => memory_space_5_sc_ack(2 downto 2),
      memory_space_5_sc_tag => memory_space_5_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 7),
      memory_space_0_lr_tag => memory_space_0_lr_tag(41 downto 21),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 16),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 7),
      memory_space_1_lr_tag => memory_space_1_lr_tag(41 downto 21),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 16),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 3),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 7),
      memory_space_2_lr_tag => memory_space_2_lr_tag(39 downto 20),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 16),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 2),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(37 downto 19),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(127 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 1),
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(1 downto 1),
      memory_space_6_lr_tag => memory_space_6_lr_tag(37 downto 19),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(31 downto 16),
      memory_space_6_lc_tag => memory_space_6_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(39 downto 20),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 16),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 2),
      memory_space_5_sr_req => memory_space_5_sr_req(1 downto 1),
      memory_space_5_sr_ack => memory_space_5_sr_ack(1 downto 1),
      memory_space_5_sr_addr => memory_space_5_sr_addr(27 downto 14),
      memory_space_5_sr_data => memory_space_5_sr_data(127 downto 64),
      memory_space_5_sr_tag => memory_space_5_sr_tag(37 downto 19),
      memory_space_5_sc_req => memory_space_5_sc_req(1 downto 1),
      memory_space_5_sc_ack => memory_space_5_sc_ack(1 downto 1),
      memory_space_5_sc_tag => memory_space_5_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(6 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(20 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(15 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(15 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(19 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(15 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(0 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(15 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(19 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(13 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(18 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(3 downto 3),
      memory_space_2_lr_ack => memory_space_2_lr_ack(3 downto 3),
      memory_space_2_lr_addr => memory_space_2_lr_addr(27 downto 21),
      memory_space_2_lr_tag => memory_space_2_lr_tag(79 downto 60),
      memory_space_2_lc_req => memory_space_2_lc_req(3 downto 3),
      memory_space_2_lc_ack => memory_space_2_lc_ack(3 downto 3),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 48),
      memory_space_2_lc_tag => memory_space_2_lc_tag(7 downto 6),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(13 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(18 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(4 downto 4),
      memory_space_0_lr_ack => memory_space_0_lr_ack(4 downto 4),
      memory_space_0_lr_addr => memory_space_0_lr_addr(34 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(104 downto 84),
      memory_space_0_lc_req => memory_space_0_lc_req(4 downto 4),
      memory_space_0_lc_ack => memory_space_0_lc_ack(4 downto 4),
      memory_space_0_lc_data => memory_space_0_lc_data(79 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(14 downto 12),
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(34 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(104 downto 84),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(79 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(14 downto 12),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(6 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(15 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(20 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(15 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(15 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(19 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(10 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(63 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(0 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(0 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(15 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(19 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_4: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 1,
      num_stores => 4,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
